// Verilog netlist created by TD v4.2.285
// Thu Dec  5 16:48:50 2019

`timescale 1ns / 1ps
module rom  // E:/WORK/RISC_V_TEST/RISC_V/al_ip/rom.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [11:0] addra;  // E:/WORK/RISC_V_TEST/RISC_V/al_ip/rom.v(18)
  input clka;  // E:/WORK/RISC_V_TEST/RISC_V/al_ip/rom.v(19)
  input rsta;  // E:/WORK/RISC_V_TEST/RISC_V/al_ip/rom.v(20)
  output [31:0] doa;  // E:/WORK/RISC_V_TEST/RISC_V/al_ip/rom.v(16)

  wire [0:1] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B0_1 ;
  wire  \inst_doa_mux_b11/B0_0 ;
  wire  \inst_doa_mux_b11/B0_1 ;
  wire  \inst_doa_mux_b12/B0_0 ;
  wire  \inst_doa_mux_b12/B0_1 ;
  wire  \inst_doa_mux_b13/B0_0 ;
  wire  \inst_doa_mux_b13/B0_1 ;
  wire  \inst_doa_mux_b14/B0_0 ;
  wire  \inst_doa_mux_b14/B0_1 ;
  wire  \inst_doa_mux_b15/B0_0 ;
  wire  \inst_doa_mux_b15/B0_1 ;
  wire  \inst_doa_mux_b16/B0_0 ;
  wire  \inst_doa_mux_b16/B0_1 ;
  wire  \inst_doa_mux_b17/B0_0 ;
  wire  \inst_doa_mux_b17/B0_1 ;
  wire  \inst_doa_mux_b18/B0_0 ;
  wire  \inst_doa_mux_b18/B0_1 ;
  wire  \inst_doa_mux_b19/B0_0 ;
  wire  \inst_doa_mux_b19/B0_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b20/B0_0 ;
  wire  \inst_doa_mux_b20/B0_1 ;
  wire  \inst_doa_mux_b21/B0_0 ;
  wire  \inst_doa_mux_b21/B0_1 ;
  wire  \inst_doa_mux_b22/B0_0 ;
  wire  \inst_doa_mux_b22/B0_1 ;
  wire  \inst_doa_mux_b23/B0_0 ;
  wire  \inst_doa_mux_b23/B0_1 ;
  wire  \inst_doa_mux_b24/B0_0 ;
  wire  \inst_doa_mux_b24/B0_1 ;
  wire  \inst_doa_mux_b25/B0_0 ;
  wire  \inst_doa_mux_b25/B0_1 ;
  wire  \inst_doa_mux_b26/B0_0 ;
  wire  \inst_doa_mux_b26/B0_1 ;
  wire  \inst_doa_mux_b27/B0_0 ;
  wire  \inst_doa_mux_b27/B0_1 ;
  wire  \inst_doa_mux_b28/B0_0 ;
  wire  \inst_doa_mux_b28/B0_1 ;
  wire  \inst_doa_mux_b29/B0_0 ;
  wire  \inst_doa_mux_b29/B0_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b30/B0_0 ;
  wire  \inst_doa_mux_b30/B0_1 ;
  wire  \inst_doa_mux_b31/B0_0 ;
  wire  \inst_doa_mux_b31/B0_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b9/B0_0 ;
  wire  \inst_doa_mux_b9/B0_1 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i0_012;
  wire inst_doa_i0_013;
  wire inst_doa_i0_014;
  wire inst_doa_i0_015;
  wire inst_doa_i0_016;
  wire inst_doa_i0_017;
  wire inst_doa_i0_018;
  wire inst_doa_i0_019;
  wire inst_doa_i0_020;
  wire inst_doa_i0_021;
  wire inst_doa_i0_022;
  wire inst_doa_i0_023;
  wire inst_doa_i0_024;
  wire inst_doa_i0_025;
  wire inst_doa_i0_026;
  wire inst_doa_i0_027;
  wire inst_doa_i0_028;
  wire inst_doa_i0_029;
  wire inst_doa_i0_030;
  wire inst_doa_i0_031;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i1_009;
  wire inst_doa_i1_010;
  wire inst_doa_i1_011;
  wire inst_doa_i1_012;
  wire inst_doa_i1_013;
  wire inst_doa_i1_014;
  wire inst_doa_i1_015;
  wire inst_doa_i1_016;
  wire inst_doa_i1_017;
  wire inst_doa_i1_018;
  wire inst_doa_i1_019;
  wire inst_doa_i1_020;
  wire inst_doa_i1_021;
  wire inst_doa_i1_022;
  wire inst_doa_i1_023;
  wire inst_doa_i1_024;
  wire inst_doa_i1_025;
  wire inst_doa_i1_026;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[10]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hCC6B6A215A683F48AA52028D94E00000054B0CF6A70000AB00000003E6666666),
    .INITP_01(256'hDAB4311C097D84F121101DAEABD6E027C053A633244D1382562368A95EBEEEEE),
    .INITP_02(256'h766D278823E42D45A8ACAE88575B74F957729F6EAF667CA0608821B8482101F6),
    .INITP_03(256'h2DC602A33320100586200A68391CAEB7FF55412A81A0303252BCE7D2A155B829),
    .INIT_00(256'h3793139313931393139313931393139313931393139313931393139313931393),
    .INIT_01(256'h1313131313131313131313131313131313131313131313736F0B232323231313),
    .INIT_02(256'h030B0393EF8B1313232323232323232323232323232323230B230B230B938B0B),
    .INIT_03(256'h00000000670B670B670B730B0B8B8303830383038303830383038303830B038B),
    .INIT_04(256'h97331313EF933313139397000000000000000000000000000000000000000000),
    .INIT_05(256'h1313131313B3B793639363939393132323239323232313231373EF139303EF93),
    .INIT_06(256'h6F33B31393EF13636703339313B76393339313333313931333B7136393639313),
    .INIT_07(256'h931333B3939313B76F93136F93E393136F33933393EF13636F13136F13E31313),
    .INIT_08(256'h6393333393B313339313333313333363B33393EF139313EF139313EF139313EF),
    .INIT_09(256'hE3136313E3139313136F1313631393133393B763931363939363936313331393),
    .INIT_0A(256'h131313376F1313E31393136313936393333333B393E313B3936F936F136F1313),
    .INIT_0B(256'h9313931323231393233323B31393131337671383038303830383331333131313),
    .INIT_0C(256'h936F1363936FB3B393139337631313631313B363136363636333936363139313),
    .INIT_0D(256'h6393B3B7E3936F9363936FB36313636333636F3333333333936F13639333B7E3),
    .INIT_0E(256'h6FE3E36F93639313631313B313376313B36363636313136FB3B3B3B3B3936F93),
    .INIT_0F(256'h33B7E313936F136393E313936F13331337E313B36313E31363636F1393B36393),
    .INIT_10(256'h6F936393B3B7E3936F939363936F93B36313636333636F13B33333333333936F),
    .INIT_11(256'h6F13B793E3E36F9393636F93B36313B3E36F936363636313136FB3B3B333B393),
    .INIT_12(256'h936F136FB33393B76F1393E36F13B3333333B3131333633313EF139333639333),
    .INIT_13(256'h6F936713830333339313139303831393B763639313B31337631313631393136F),
    .INIT_14(256'h231367136F33339367336333136393336733133763936393B393139313376F93),
    .INIT_15(256'h136313671383038333331313939313331363136313B393EF1393333393632323),
    .INIT_16(256'h6F9393136F13B3933393B7639313639313633393133733136313333333339333),
    .INIT_17(256'h93B3B33333B3B3136393333313B7639363639393631393939333131393131313),
    .INIT_18(256'h936FB71363936FB363B36FB333931333136FB3B3B3B3136393B393B3936F6313),
    .INIT_19(256'h6F936F93E3131393936733B3939393939393B763639313B31337631393631393),
    .INIT_1A(256'h13EF9367E3139333B36313E3931363639363139313636367E313933363931313),
    .INIT_1B(256'h1337B3331393B39363B76733EF33E3B36713EF6363936733EF93B36FB3633367),
    .INIT_1C(256'h6F93A393938363939367E3A393938363936393633393B36F93E39337673303B3),
    .INIT_1D(256'h1367E3E3239393036F2393232323232323230323938303038303838383631393),
    .INIT_1E(256'h23A323A323A323A323A32367B39793B36763E31323232323B313936363936313),
    .INIT_1F(256'h132313671333E30393936FE333339393E793B397936FB393B393936723A323A3),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n63,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_008,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0290C09080FE2C02600000004220000000000000000000000000000000000000),
    .INITP_01(256'hA0427F3E6DDBF73AA33F654513E1FC54C152000301128558AA085244AEFDEC84),
    .INITP_02(256'h3A92494A8EDC48A1400C54100A2D40B2C0505619F28A400D0C6FBCCEA8A5F795),
    .INITP_03(256'h07BFAC0FFFFB7FEE3AFFD007EA3455075628A2914E1D4048BA379DAE5A766453),
    .INIT_00(256'h2007070707060606060505050504040404030303030202020201010101000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000030939291908080),
    .INIT_02(256'h509050800862020057565554515057565554535257565552E051A05020009050),
    .INIT_03(256'h00000000406240B240B20000A060575757575454535353535252515151905090),
    .INIT_04(256'h120303020002030302C000000000000000000000000000000000000000000000),
    .INIT_05(256'hBA4A6A058472034A810383AC6AC5BC9296978A919395AC9480000803829200C2),
    .INIT_06(256'hF8844A0483004245809383438B137784E4038384B30B038232030A8403866D2A),
    .INIT_07(256'h02423A7A2B6F4787F80302F803000302F8C2030A83000205F80504F805430504),
    .INIT_08(256'hEE0BF233CBC3AB1AEB8A83B98BFB82FAC383AB00C2C28700C202830042C28100),
    .INIT_09(256'hCC03C703C1030342C4000302EC2A03433AC303ED0B02C2033BC53B2B43F23A2B),
    .INIT_0A(256'h0A040302000302E92A0B02C2033BC53BF21A0A2B44A603C303F884F844000302),
    .INIT_0B(256'hCB44AA0392933C7B90BB91BBECAB838003408095959494929290320A322A8BBB),
    .INIT_0C(256'h0200024F0200F3FBEB83FB03870382AECB42C30F03830E2ECF43E28A0A8BEA02),
    .INIT_0D(256'h6B03F3030503F8830F03F8C30B03C64A0303F8B31B8BC3AA02F803EB02B30245),
    .INIT_0E(256'h0087C300C38103FB84FB02FB8303ADCBC380C2498D3A43F8F31BCBEA4303F803),
    .INIT_0F(256'hB3024102020003E9024002020084FA0202A8CBC3090385420C2CF802EBC30003),
    .INIT_10(256'hF8036B03F3030403F8C2830803F8C2830C03C04C0305F842C3B31B8BC3AA02F8),
    .INIT_11(256'h000203028ACC00020348F8C2832C4BC387008383CC488FBA42F8331BCBEC4303),
    .INIT_12(256'h83F842F83B82C303F8020309F802F31A0A822B038282A70A820002C2826A0BC2),
    .INIT_13(256'hF84340809294B2B24AEA8BCB9290BA0203C38CEB03FB8303810382AFCB0302F8),
    .INIT_14(256'h93804002F8AAC3034002408A83EE03F24042A202FD02FBABFB02BB03AB03F803),
    .INIT_15(256'h03A803408092929032324A2ACBFB0A0A82AB03A103C3030002AA02E2AB829192),
    .INIT_16(256'hF8020302F8AAC303BBC3036E8B8302033A453B3B83030A83AB03B21A0A2B8383),
    .INIT_17(256'h03B3F3AA0B1B8B04E40382330203660320E10303C38BEAFB0333AB3C0BEC2BCB),
    .INIT_18(256'h03F8030BC603F81B0B33F833B3AB0B1A8AF8731B730C0483042B03C3030080FB),
    .INIT_19(256'hF803F8C38603FB030340F2F3CAEB4B7BCB0203C34CEB03FB8303410343AFCB03),
    .INIT_1A(256'hC2F841404B2B6BB2C2F302354B0B2C3D03060282C3E3A040CB0BEA8242FB0283),
    .INIT_1B(256'h8212AB8303CBDB03BD834002F802AC0240C2F8A6E5414002F84102F802EC0240),
    .INIT_1C(256'hF8FBC7C2C3E34783BB40F4C7C2C3E3BE83F103CB83FBE3F803B503034082E2C3),
    .INIT_1D(256'h0140F4F4D7C2C3D3F8D7C3D7D6D5D4D3D2D1D4D0C2D4D1D7D7D7D7D1D1FA43BB),
    .INIT_1E(256'h81818181828282828383834043014B83400AB38393929190433B3BC9C8BBBF83),
    .INIT_1F(256'h8293804082C28EE3C383F8BC0383C34040414301CBF8F2CBF2CBFA4080808080),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n106,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_017,inst_doa_i0_016,inst_doa_i0_015,inst_doa_i0_014,inst_doa_i0_013,inst_doa_i0_012,inst_doa_i0_011,inst_doa_i0_010,inst_doa_i0_009}));
  // address_offset=0;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h029588958C00204882420081002000000053F00000FC00000000004200000000),
    .INITP_01(256'h783984A1E00C3C021C644003EC540E8013030001200004542822400800001110),
    .INITP_02(256'h0001611088600D00000490044808227080020BC3531000C448000700870C4401),
    .INITP_03(256'h2B1204200000202038402007A0300140810A200008102680000102F14400400C),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h000000000000000000000000000000000000000000000004E08000000000C000),
    .INIT_02(256'h1080000120000000FCF8F4F04440BCB8B4B0ACA81C1814080008000800008080),
    .INIT_03(256'h0000000000000081008104000000F0E0D0C01000F0E0D0C0B0A0706050802080),
    .INIT_04(256'h002920004400294020B0FF000000000000000000000000000000000000000000),
    .INIT_05(256'hFD265E00063D000DBEFC027D2501FE50200425544C245D488004100010008471),
    .INIT_06(256'hD72A3D28EDC4018101013571090039065638FD2A3D0A00053D000DBDFC017E25),
    .INIT_07(256'h010171714141FF00370400670C8108FCA729283DEDC40181670400970C8108FC),
    .INIT_08(256'h011139391929692041191970417175793979404403010184030101C401010104),
    .INIT_09(256'h3904B90CB90802010290FC00B90DF8023DFD0001111135103D011D38FE210505),
    .INIT_0A(256'h2500FC10400400810D151139103D011D2120453D7A3D6C3904D7026702D00000),
    .INIT_0B(256'h0D017DFC2004FEFD482D24295D5DFDC020008010203040506070297E39255DFD),
    .INIT_0C(256'hFC80FC2DFCC0353905FD0580B9FC050115013981FD010230A5410501320D7D02),
    .INIT_0D(256'h316C3500B6FC470136FCA73901FD81813681073938313131807704316C2D00AD),
    .INIT_0E(256'hD081817011B5103D811D0439FD0001153981010101F905C73D3C353131803704),
    .INIT_0F(256'h2D00ADFCFCD004B16C2DFCFC200121FD0081153981FD810102301701053935FC),
    .INIT_10(256'h1704316C3500B6FC670101B6FCB7013D01FD0181368147013939383131318077),
    .INIT_11(256'h40FC80008101A000008117013D01153901600181010101F905A73E3C35313180),
    .INIT_12(256'h018701A73D2AFD001700000137002120292929800549C929ED0001013D011539),
    .INIT_13(256'h77010040100025397D255D252030FD001001390DFC39FD00B9FC05011500FC67),
    .INIT_14(256'h04C00000A739395800288139A93954310029FD003974397D29F8FDFD5D20A700),
    .INIT_15(256'h14BD640040102030293D7D255DFD2529E129203D582978E0017D3D297D812420),
    .INIT_16(256'h27000000670D297C3DFD0001151135103D01391DFD0039ED2914212035396D29),
    .INIT_17(256'h003D3129413C410AA97C353D78203DA43435F802810D7DF9063D75FE0D513131),
    .INIT_18(256'h0067800D01FC673C0239B73D31750D2819173D3C3A418A3D00358035F870011D),
    .INIT_19(256'hA700471131103D0004002D357D255DFD25001001390DFC39FD00B9FC050115FC),
    .INIT_1A(256'h01D7000081050535313100AD0505302D0481FC01018181008105053101050001),
    .INIT_1B(256'h61003D3D800D29FCBD00002C8728812C0001E7010100002847002C772C012800),
    .INIT_1C(256'hA70DB505050101010D00B9B5050501B901B10C01310D29376039404000290129),
    .INIT_1D(256'h3C0039B5B1111101B7C19145197175797D15F11D917161514131211101B181F1),
    .INIT_1E(256'h2D2D2D2D2D2D2D2D2D2D2D31150009300001B5412D2D2D2D393DC101813DB001),
    .INIT_1F(256'hC0A04000FD2981FD0501F7B03D3DC1008100150009B735413521FD002D2D2D2D),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n149,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_026,inst_doa_i0_025,inst_doa_i0_024,inst_doa_i0_023,inst_doa_i0_022,inst_doa_i0_021,inst_doa_i0_020,inst_doa_i0_019,inst_doa_i0_018}));
  // address_offset=0;data_offset=27;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00010000000000000081000000000000000000000000C00C0000000000000000),
    .INIT_01(256'h000C82218CC0822183C000040C03015040C054040000C40D04417C0000000000),
    .INIT_02(256'h0105000F000000010403000000702300C0C014453C0001004000000001010102),
    .INIT_03(256'h09403583303C1C01980000F00013000C00DC18340C0030035450339200E18000),
    .INIT_04(256'h80000004004F1007330FC3000000D0005094240040013000C00D0060340C0003),
    .INIT_05(256'h0001000B5543030080813C0000F3000004000010C046001030C100840C10070C),
    .INIT_06(256'h0001008C0800C30030C003000C00C000CCC000010004F101301C0C00300400D4),
    .INIT_07(256'h0CCF0A0CC0200400000000000C000D400BC0F0000C00000FCC000F0100033000),
    .INIT_08(256'h0C03F2010FDFFFCC3CCFFC030033C333030030C0C00FFF0CCCF0300FF00CCCFF),
    .INIT_09(256'h0300C00333FFCCCE0F8FFF30F33FC0330030043C83202C3F3FFF03000EFF44F2),
    .INIT_0A(256'hC03336FF84C84C3CC310FCC083F7F3FF00F33FCCFCFC7CCC04033CD00037CF00),
    .INIT_0B(256'hD1173CC4F040CF0F30523D1DDF403000E3CF3C333033303304CCCCF7CCCCFC3C),
    .INIT_0C(256'h00CC03302CC07300C80345010CC51C00D803A00E803A00FC0EE0FCD1E0031315),
    .INIT_0D(256'h0A0A0A0E0E0A0A0A0A0A0A0A111F068540000000000000E000FC00FC00FC003F),
    .INIT_0E(256'h0000000000000000000005555555555555555000000000000000000000000A0A),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_027 (
    .addra({addra,1'b1}),
    .clka(clka),
    .dia({open_n198,open_n199,open_n200,1'b0,open_n201,open_n202,1'b0,open_n203,open_n204}),
    .rsta(rsta),
    .doa({open_n219,open_n220,open_n221,open_n222,open_n223,open_n224,open_n225,inst_doa_i0_028,inst_doa_i0_027}));
  // address_offset=0;data_offset=29;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000C1000000000000000000000000000C0000000000000000),
    .INIT_01(256'h000CC330ECD0C330E3D002000C03000000C000000000C80524896C0000000000),
    .INIT_02(256'h0000000F000000000003000000323300C0C000003C0000000000000000000000),
    .INIT_03(256'h0C003003323C0C043D1040F00403008C00CC0C348C0830030000334000D02000),
    .INIT_04(256'h80000000000F0002222FC3C02020E08200F00C82C0003008C00CC032308C8083),
    .INIT_05(256'h0002080302030300C0C83C0000F3000200000000C021088030C820C00C00030C),
    .INIT_06(256'h820002EE0C02CB8830C083000C00C000CCC000000000F000300C0C00300802C0),
    .INIT_07(256'h0CEF0F2CC0300000000000020C000C000FC0F0000C00000FCC000F0000033020),
    .INIT_08(256'h0CC3F1030FCFFFC43CCFFC030033C333030030C0C00FFF2CCCF0300FF00CCCFF),
    .INIT_09(256'h0300C00333EFECCE0F8EFF00F33FC4330430043CC3101C3F3FFF03000FFFC0F1),
    .INIT_0A(256'h803333FF40C40C3CC310FCC043F3F3FF82F33FCCCCFCBCCC04133CD40437CF00),
    .INIT_0B(256'hD1173CC0F202CF1720593D2D13403000E3CF30333433343340CCCC37CCCCFCBC),
    .INIT_0C(256'h02F407D00F403D00F40345010CC51C00F403D00F403D00FC0FD0FCD150031315),
    .INIT_0D(256'hC7C7C7C7C7C7C7C7C7C7C7C7E007C3C3C0000000000000E800E400E400E40039),
    .INIT_0E(256'h00000000000000000000000000000000000000000000000000000000000007C7),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_029 (
    .addra({addra,1'b1}),
    .clka(clka),
    .dia({open_n257,open_n258,open_n259,1'b0,open_n260,open_n261,1'b0,open_n262,open_n263}),
    .rsta(rsta),
    .doa({open_n278,open_n279,open_n280,open_n281,open_n282,open_n283,open_n284,inst_doa_i0_030,inst_doa_i0_029}));
  // address_offset=0;data_offset=31;depth=4096;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000040000000000000000),
    .INIT_01(256'h0004411044404110414001000401000000400000000040010000140000000000),
    .INIT_02(256'h0000000500000000000100000010110040400000140000000000000000000000),
    .INIT_03(256'h0400100110140400140000500001000400440410040010010000100000400000),
    .INIT_04(256'h4000000000050001110541400000400000500400400010004004401010040001),
    .INIT_05(256'h0001000101000000404014000051000000000000400000001040004005000104),
    .INIT_06(256'h4000004404004100104001000400400044400000000050001004040010040040),
    .INIT_07(256'h0445050440100000000000000400040005405000040000054400050000011000),
    .INIT_08(256'h0441510105455544144554010011411101001040400555144450100550044455),
    .INIT_09(256'h0100400111554445054555105115441104100414411014151555010005554051),
    .INIT_0A(256'h4011115540440414411054404151515500511544445454440401144000114500),
    .INIT_0B(256'h4001144050004511100515140140100051451411141114114044445544445454),
    .INIT_0C(256'h0054015005401500540100000440040054015005401500540550544050010100),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000540054005400540115),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_031 (
    .addra({addra,1'b1}),
    .clka(clka),
    .dia({open_n316,open_n317,open_n318,open_n319,open_n320,open_n321,1'b0,open_n322,open_n323}),
    .rsta(rsta),
    .doa({open_n338,open_n339,open_n340,open_n341,open_n342,open_n343,open_n344,open_n345,inst_doa_i0_031}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00A7F2F684ABB15CDDDD6FBAA0146B7AF7EEF155D901436C147CA66B9056DD9C),
    .INITP_01(256'h74DBDF8ABDCAAC51B6DCDCD3767559F573CF79ED7BF778BAFF559F56FBD95CC0),
    .INITP_02(256'h00000000000014B88000109BBBBBBBBDDBB76EDDBB6B6F7DBB76EDD8275B777C),
    .INITP_03(256'h00C000000000000000000000000000000000000000000000003FFFC03CE2B200),
    .INIT_00(256'h836F23932323132323136713031383E383032393B7032313836F23B383032323),
    .INIT_01(256'h1323231367130313230393B7A393132313671303831383E32313832393EF0393),
    .INIT_02(256'h93832393836F238323232313232323136713038313E38383EF13832313836F23),
    .INIT_03(256'h13938313EF13939383A393EF139393EF13939383836F23832383E3832393EF13),
    .INIT_04(256'h93EF0323232323231323231367138303831383E383239383EF139393832393EF),
    .INIT_05(256'h9393EF13938363931393EF1393832393EF1393EF1383B71393EF039393EF0323),
    .INIT_06(256'h136F2323EF1323EF03E3832393EF1393832393836F2323832393EF1393836F23),
    .INIT_07(256'h2323232313232323136713038313B3833383138323EF03E303B38313239383EF),
    .INIT_08(256'h83B393B71363139383832393836F63136313631383836F239393232323232323),
    .INIT_09(256'h93B3131383A393836FA3238323832313836F23B30383A393EF03238323138367),
    .INIT_0A(256'hEF13938313EF13939383A393EF139393EF13939383836F238323B30383E38323),
    .INIT_0B(256'hEF9313830323139393836FE383A39383EF139393836FEF139393836393032393),
    .INIT_0C(256'hEF1393832313836F23B38313EF03EF0323832313836F23B30383A393EF032393),
    .INIT_0D(256'h83E38383239383239383EF1383836F239383EF1383836F239383EF1313239383),
    .INIT_0E(256'h93EF13938303EF13B78323EF13EF03231323132393B713232313671383038313),
    .INIT_0F(256'hEF139383638323E3B7032393832313B3038393B313339393036F2323B7EF1323),
    .INIT_10(256'h2323136FEF13B793E383239383231383EF13B7931383B3839383338313832323),
    .INIT_11(256'h83EF13B793639383EF13B793639383EF13B793639383EF13B793639383232313),
    .INIT_12(256'h83EF13B79363938323138323136393036393032303B393036383A38393B76393),
    .INIT_13(256'hB793639383EF13B793639383EF13B793639383EF13B793639383EF13B7936393),
    .INIT_14(256'h9363B3B703EF13B79363B3B703EF13B79363B3B703EF13B79363B393B703EF13),
    .INIT_15(256'h68BC909090902C909090909090909090909090D8908464671303831383EF13B7),
    .INIT_16(256'h490D7472490D7472490D7472490D74724980007A0A202572200A3D6B200A726F),
    .INIT_17(256'h490D7472490D7472490D7472490D7472490D7472490D7472490D7472490D7472),
    .INIT_18(256'h0606050505050404030070DCDCDC0CE070E00C70E0E00CE8E80D7472490D7472),
    .INIT_19(256'h0808080808080808080807070707070707070707070707070707060606060606),
    .INIT_1A(256'h0000000000000000000008080808080808080808080808080808080808080808),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000D0E800000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n371,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_008,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=1024;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0006A54509462030B2B0DF54400052F1CB156023100006E800A0054500053510),
    .INITP_01(256'hA9173F0473940C0164B8B8A2F44A5108BB92F3D0E58AB024F2051095FD92A880),
    .INITP_02(256'h00000000000000117FFFFE1767676773B76EDDBB7644949B76EDDBB01E92FEA8),
    .INITP_03(256'h000000000000000000000000000000000000000000000000003FFFFFC0FFFF80),
    .INIT_00(256'h13001303161782929380408092C2138F1313D0C303E317C31300138313131617),
    .INIT_01(256'h8296978040809200D023C303038382978040809290C213CF16C3131383F812C2),
    .INIT_02(256'h021313C31300121311131782919293804080929000C8E313F8C2E313C3130013),
    .INIT_03(256'hC2821383F802C2C3130083F842C283F802C2C313120012131113CE131283F8C2),
    .INIT_04(256'h83F8121213161713829697804080929290C213CF1313C313F8C2FBC3231283F8),
    .INIT_05(256'hC383F8C20213E903C383F8C202131183F8C283F082D213C383F812C283F81215),
    .INIT_06(256'h02001010F80217F812CE131283F8C2021313C313001312131183F8C202130011),
    .INIT_07(256'h13121113829596978040809290C283138313C31316F812A71383130310C313F8),
    .INIT_08(256'hD383C313CBB203C3E31313C31300C303C403C503E3130014C303111017161514),
    .INIT_09(256'hEB83BBEB1302C3230002131317D314C31300118313230283F81217D314C313C0),
    .INIT_0A(256'hF8C2821383F802C2C3230683F842C283F802C2C3231200131311831323CE1313),
    .INIT_0B(256'hF802C2D3D414C3FBC31300CE2302C323F8C2FBC32300F8C2FBC323F703231383),
    .INIT_0C(256'hF8C2FBD314C3130011831383F812F81210D314C31300118313230283F8121583),
    .INIT_0D(256'h13CCE31313C31311C313F8C2E3130011C313F8C2E3130011C313F8020011C313),
    .INIT_0E(256'h83F882C21313F8C2131210F002F8121103100311C313829293804080929290C2),
    .INIT_0F(256'hF802C213C01310A7231312C313C07B831313C383BB83EBAB1300121703F00213),
    .INIT_10(256'h929380F8F8C21302CB1313C31310C313F8C21382C3E3C313C313C313C3131312),
    .INIT_11(256'h13F8C21302C5FB13F8C21302C5FB13F8C21302C5FB13F8C21302C5FB13161782),
    .INIT_12(256'h13F8C21302C5FB1312C3131303FB0313840323C023830313C91303E3C303C7FB),
    .INIT_13(256'h1302C5FB13F8C21302C5FB13F8C21302C5FB13F8C21302C5FB13F8C21302C5FB),
    .INIT_14(256'h02C5BB2313F8C21302C5BB1313F8C21302C5BB0B13F8C21302C5BBC30B13F8C2),
    .INIT_15(256'h320A0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0A0B0A0B40809290C213F8C213),
    .INIT_16(256'h370510B9370510B9370510B9370510B9374B001E00123C1030001234B6003690),
    .INIT_17(256'h370590B9370590B9370590B9370510B9370510B9370510B9370510B9370510B9),
    .INIT_18(256'h030382828282020281000202020202020202020202020202020590B9370590B9),
    .INIT_19(256'h0404040404040404040483838383838383838383838383838383030303030303),
    .INIT_1A(256'h0000000000000000000004040404040404040404040404040404040404040404),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000030100000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_001024_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n414,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_017,inst_doa_i1_016,inst_doa_i1_015,inst_doa_i1_014,inst_doa_i1_013,inst_doa_i1_012,inst_doa_i1_011,inst_doa_i1_010,inst_doa_i1_009}));
  // address_offset=1024;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h18215BAA3BF4D785042690273F903F2D29D03BF86BE10515104883F6AC43C2AF),
    .INITP_01(256'h886AC8F70262BB909B654745AAA5AEEE055F38A694E81DDF0D7AEE6A006A27B0),
    .INITP_02(256'h88888AAA888884A38000000C0A0A0E0708103061E10228A2E142860E30680110),
    .INITP_03(256'h000000000000000000000000000000000000000000000000003FFFFFFF000028),
    .INIT_00(256'h7170BD042D29C0A0844000C0B001613DB1713921800139057180BD3D61712D29),
    .INIT_01(256'h802004800080700039BD2180BD0180208000C0A0B001B10139FD61BD01E7B101),
    .INIT_02(256'h28A1BD05B1A0BD71818129C0A4A0844000806070008101B1870101B905B170A9),
    .INIT_03(256'h0101A101B72801FDB1BD0177010101672801FDB1A110BD71BDB101A1BD018701),
    .INIT_04(256'h014331818101012900A0840000C090A0B0019181B1BDFDB18701FDC18DBD01D7),
    .INIT_05(256'h0501C7012891B910010157012891BD01330101B701E100010193310101C3513D),
    .INIT_06(256'hC060818147B829875101A1BD01770128A1BD05B1A081BD91BD014701289170BD),
    .INIT_07(256'h35312D2900A4A084800000E0F0013D613DB105712967913D813DB118BD0581F7),
    .INIT_08(256'h013D910009BD547501313D05310039283994B9340131303D9181818145413D39),
    .INIT_09(256'h113D3D7DB1BD05ADA081BD713D0139114160BD3D91ADBD0197713D0139114101),
    .INIT_0A(256'hE30101B101C74001FDAD3D0183010101774001FDADB1A0BD71BD3D91AD01B1BD),
    .INIT_0B(256'h13020101113921E11D41F001ADBDFDAD0701FD5D6D606701FDC16D39246DBD01),
    .INIT_0C(256'h0701FD01391141C0BD3D91013781B781BD01391141A0BD3D91ADBD0117513D01),
    .INIT_0D(256'h918101313D0531BD0591A701013180BD05912701013100BD0591A72800BD0591),
    .INIT_0E(256'h012301011000E7310081A92700579138D038D0BDF100402004C00080D0E0F001),
    .INIT_0F(256'hE3400120813000BD00A1BD05A139FD3D71A1013DFD3D617DA100813DC067A0BD),
    .INIT_10(256'hA08440E723C1001001B1BD05B138050087710001010135710100397101000000),
    .INIT_11(256'h61F3B1003801216163710038011161D331003801096143F100380105612D29C0),
    .INIT_12(256'h61F3F100380181613805203804398C203D28BD39BD3D40200130BD0121800141),
    .INIT_13(256'h003801016133F10038010161A3B1003801016113710038010161833100380101),
    .INIT_14(256'h38013D006133F10038013D0061B3B10038013D006133710038013D010061C331),
    .INIT_15(256'h1B0000000000000000000000000000000000000000000000C0A0B00171B33100),
    .INIT_16(256'h5D00C81D5D00881D5D00481D5D00081D5DC6008C005E880C19005E5CD80059DD),
    .INIT_17(256'h5D008C1D5D004C1D5D000C1D5D00481D5D00081D5D00C81D5D00881D5D00481D),
    .INIT_18(256'h8181414141410101C080000000000000000000000000000000000C1D5D00CC1D),
    .INIT_19(256'h02020202020202020202C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1818181818181),
    .INIT_1A(256'h0000000000000000000002020202020202020202020202020202020202020202),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_001024_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n457,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_026,inst_doa_i1_025,inst_doa_i1_024,inst_doa_i1_023,inst_doa_i1_022,inst_doa_i1_021,inst_doa_i1_020,inst_doa_i1_019,inst_doa_i1_018}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n500,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_008,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n543,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_008,inst_doa_i3_007,inst_doa_i3_006,inst_doa_i3_005,inst_doa_i3_004,inst_doa_i3_003,inst_doa_i3_002,inst_doa_i3_001,inst_doa_i3_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i1_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b10/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i1_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b11/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_0  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i1_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b12/B0_0 ),
    .i1(\inst_doa_mux_b12/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[12]));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_0  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i1_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b13/B0_0 ),
    .i1(\inst_doa_mux_b13/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[13]));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_0  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i1_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b14/B0_0 ),
    .i1(\inst_doa_mux_b14/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[14]));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_0  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i1_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b15/B0_0 ),
    .i1(\inst_doa_mux_b15/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[15]));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_0  (
    .i0(inst_doa_i0_016),
    .i1(inst_doa_i1_016),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_0 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_1 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b16/B0_0 ),
    .i1(\inst_doa_mux_b16/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[16]));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_0  (
    .i0(inst_doa_i0_017),
    .i1(inst_doa_i1_017),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_0 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_1 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b17/B0_0 ),
    .i1(\inst_doa_mux_b17/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[17]));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_0  (
    .i0(inst_doa_i0_018),
    .i1(inst_doa_i1_018),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_0 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_1 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b18/B0_0 ),
    .i1(\inst_doa_mux_b18/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[18]));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_0  (
    .i0(inst_doa_i0_019),
    .i1(inst_doa_i1_019),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_0 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_1 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b19/B0_0 ),
    .i1(\inst_doa_mux_b19/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[19]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_0  (
    .i0(inst_doa_i0_020),
    .i1(inst_doa_i1_020),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_0 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_1 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b20/B0_0 ),
    .i1(\inst_doa_mux_b20/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[20]));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_0  (
    .i0(inst_doa_i0_021),
    .i1(inst_doa_i1_021),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_0 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_1 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b21/B0_0 ),
    .i1(\inst_doa_mux_b21/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[21]));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_0  (
    .i0(inst_doa_i0_022),
    .i1(inst_doa_i1_022),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_0 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_1 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b22/B0_0 ),
    .i1(\inst_doa_mux_b22/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[22]));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_0  (
    .i0(inst_doa_i0_023),
    .i1(inst_doa_i1_023),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_0 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_1 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b23/B0_0 ),
    .i1(\inst_doa_mux_b23/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[23]));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_0  (
    .i0(inst_doa_i0_024),
    .i1(inst_doa_i1_024),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_0 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_1 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b24/B0_0 ),
    .i1(\inst_doa_mux_b24/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[24]));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_0  (
    .i0(inst_doa_i0_025),
    .i1(inst_doa_i1_025),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_0 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_1 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b25/B0_0 ),
    .i1(\inst_doa_mux_b25/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[25]));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_0  (
    .i0(inst_doa_i0_026),
    .i1(inst_doa_i1_026),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_0 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_1 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b26/B0_0 ),
    .i1(\inst_doa_mux_b26/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[26]));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_0  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_0 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_1  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_1 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b27/B0_0 ),
    .i1(\inst_doa_mux_b27/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[27]));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_0  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_0 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_1  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_1 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b28/B0_0 ),
    .i1(\inst_doa_mux_b28/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[28]));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_0  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_0 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_1  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_1 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b29/B0_0 ),
    .i1(\inst_doa_mux_b29/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[29]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_0  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_0 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_1  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_1 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b30/B0_0 ),
    .i1(\inst_doa_mux_b30/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[30]));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_0  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_0 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_1  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_1 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b31/B0_0 ),
    .i1(\inst_doa_mux_b31/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[31]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i1_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b9/B0_0 ),
    .i1(\inst_doa_mux_b9/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[9]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

