// Verilog netlist created by TD v4.2.285
// Wed Jun 17 17:40:49 2020

`timescale 1ns / 1ps
module rom  // E:/WORK/RISC_V_TEST/picorv32_EG4S20/RISC_V/al_ip/rom.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [12:0] addra;  // E:/WORK/RISC_V_TEST/picorv32_EG4S20/RISC_V/al_ip/rom.v(18)
  input clka;  // E:/WORK/RISC_V_TEST/picorv32_EG4S20/RISC_V/al_ip/rom.v(19)
  input rsta;  // E:/WORK/RISC_V_TEST/picorv32_EG4S20/RISC_V/al_ip/rom.v(20)
  output [31:0] doa;  // E:/WORK/RISC_V_TEST/picorv32_EG4S20/RISC_V/al_ip/rom.v(16)

  wire [0:2] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B0_2 ;
  wire  \inst_doa_mux_b0/B0_3 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b0/B1_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B0_2 ;
  wire  \inst_doa_mux_b1/B0_3 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b1/B1_1 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B0_1 ;
  wire  \inst_doa_mux_b10/B0_2 ;
  wire  \inst_doa_mux_b10/B0_3 ;
  wire  \inst_doa_mux_b10/B1_0 ;
  wire  \inst_doa_mux_b10/B1_1 ;
  wire  \inst_doa_mux_b11/B0_0 ;
  wire  \inst_doa_mux_b11/B0_1 ;
  wire  \inst_doa_mux_b11/B0_2 ;
  wire  \inst_doa_mux_b11/B0_3 ;
  wire  \inst_doa_mux_b11/B1_0 ;
  wire  \inst_doa_mux_b11/B1_1 ;
  wire  \inst_doa_mux_b12/B0_0 ;
  wire  \inst_doa_mux_b12/B0_1 ;
  wire  \inst_doa_mux_b12/B0_2 ;
  wire  \inst_doa_mux_b12/B0_3 ;
  wire  \inst_doa_mux_b12/B1_0 ;
  wire  \inst_doa_mux_b12/B1_1 ;
  wire  \inst_doa_mux_b13/B0_0 ;
  wire  \inst_doa_mux_b13/B0_1 ;
  wire  \inst_doa_mux_b13/B0_2 ;
  wire  \inst_doa_mux_b13/B0_3 ;
  wire  \inst_doa_mux_b13/B1_0 ;
  wire  \inst_doa_mux_b13/B1_1 ;
  wire  \inst_doa_mux_b14/B0_0 ;
  wire  \inst_doa_mux_b14/B0_1 ;
  wire  \inst_doa_mux_b14/B0_2 ;
  wire  \inst_doa_mux_b14/B0_3 ;
  wire  \inst_doa_mux_b14/B1_0 ;
  wire  \inst_doa_mux_b14/B1_1 ;
  wire  \inst_doa_mux_b15/B0_0 ;
  wire  \inst_doa_mux_b15/B0_1 ;
  wire  \inst_doa_mux_b15/B0_2 ;
  wire  \inst_doa_mux_b15/B0_3 ;
  wire  \inst_doa_mux_b15/B1_0 ;
  wire  \inst_doa_mux_b15/B1_1 ;
  wire  \inst_doa_mux_b16/B0_0 ;
  wire  \inst_doa_mux_b16/B0_1 ;
  wire  \inst_doa_mux_b16/B0_2 ;
  wire  \inst_doa_mux_b16/B0_3 ;
  wire  \inst_doa_mux_b16/B1_0 ;
  wire  \inst_doa_mux_b16/B1_1 ;
  wire  \inst_doa_mux_b17/B0_0 ;
  wire  \inst_doa_mux_b17/B0_1 ;
  wire  \inst_doa_mux_b17/B0_2 ;
  wire  \inst_doa_mux_b17/B0_3 ;
  wire  \inst_doa_mux_b17/B1_0 ;
  wire  \inst_doa_mux_b17/B1_1 ;
  wire  \inst_doa_mux_b18/B0_0 ;
  wire  \inst_doa_mux_b18/B0_1 ;
  wire  \inst_doa_mux_b18/B0_2 ;
  wire  \inst_doa_mux_b18/B0_3 ;
  wire  \inst_doa_mux_b18/B1_0 ;
  wire  \inst_doa_mux_b18/B1_1 ;
  wire  \inst_doa_mux_b19/B0_0 ;
  wire  \inst_doa_mux_b19/B0_1 ;
  wire  \inst_doa_mux_b19/B0_2 ;
  wire  \inst_doa_mux_b19/B0_3 ;
  wire  \inst_doa_mux_b19/B1_0 ;
  wire  \inst_doa_mux_b19/B1_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b2/B0_2 ;
  wire  \inst_doa_mux_b2/B0_3 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b2/B1_1 ;
  wire  \inst_doa_mux_b20/B0_0 ;
  wire  \inst_doa_mux_b20/B0_1 ;
  wire  \inst_doa_mux_b20/B0_2 ;
  wire  \inst_doa_mux_b20/B0_3 ;
  wire  \inst_doa_mux_b20/B1_0 ;
  wire  \inst_doa_mux_b20/B1_1 ;
  wire  \inst_doa_mux_b21/B0_0 ;
  wire  \inst_doa_mux_b21/B0_1 ;
  wire  \inst_doa_mux_b21/B0_2 ;
  wire  \inst_doa_mux_b21/B0_3 ;
  wire  \inst_doa_mux_b21/B1_0 ;
  wire  \inst_doa_mux_b21/B1_1 ;
  wire  \inst_doa_mux_b22/B0_0 ;
  wire  \inst_doa_mux_b22/B0_1 ;
  wire  \inst_doa_mux_b22/B0_2 ;
  wire  \inst_doa_mux_b22/B0_3 ;
  wire  \inst_doa_mux_b22/B1_0 ;
  wire  \inst_doa_mux_b22/B1_1 ;
  wire  \inst_doa_mux_b23/B0_0 ;
  wire  \inst_doa_mux_b23/B0_1 ;
  wire  \inst_doa_mux_b23/B0_2 ;
  wire  \inst_doa_mux_b23/B0_3 ;
  wire  \inst_doa_mux_b23/B1_0 ;
  wire  \inst_doa_mux_b23/B1_1 ;
  wire  \inst_doa_mux_b24/B0_0 ;
  wire  \inst_doa_mux_b24/B0_1 ;
  wire  \inst_doa_mux_b24/B0_2 ;
  wire  \inst_doa_mux_b24/B0_3 ;
  wire  \inst_doa_mux_b24/B1_0 ;
  wire  \inst_doa_mux_b24/B1_1 ;
  wire  \inst_doa_mux_b25/B0_0 ;
  wire  \inst_doa_mux_b25/B0_1 ;
  wire  \inst_doa_mux_b25/B0_2 ;
  wire  \inst_doa_mux_b25/B0_3 ;
  wire  \inst_doa_mux_b25/B1_0 ;
  wire  \inst_doa_mux_b25/B1_1 ;
  wire  \inst_doa_mux_b26/B0_0 ;
  wire  \inst_doa_mux_b26/B0_1 ;
  wire  \inst_doa_mux_b26/B0_2 ;
  wire  \inst_doa_mux_b26/B0_3 ;
  wire  \inst_doa_mux_b26/B1_0 ;
  wire  \inst_doa_mux_b26/B1_1 ;
  wire  \inst_doa_mux_b27/B0_0 ;
  wire  \inst_doa_mux_b27/B0_1 ;
  wire  \inst_doa_mux_b27/B0_2 ;
  wire  \inst_doa_mux_b27/B0_3 ;
  wire  \inst_doa_mux_b27/B1_0 ;
  wire  \inst_doa_mux_b27/B1_1 ;
  wire  \inst_doa_mux_b28/B0_0 ;
  wire  \inst_doa_mux_b28/B0_1 ;
  wire  \inst_doa_mux_b28/B0_2 ;
  wire  \inst_doa_mux_b28/B0_3 ;
  wire  \inst_doa_mux_b28/B1_0 ;
  wire  \inst_doa_mux_b28/B1_1 ;
  wire  \inst_doa_mux_b29/B0_0 ;
  wire  \inst_doa_mux_b29/B0_1 ;
  wire  \inst_doa_mux_b29/B0_2 ;
  wire  \inst_doa_mux_b29/B0_3 ;
  wire  \inst_doa_mux_b29/B1_0 ;
  wire  \inst_doa_mux_b29/B1_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b3/B0_2 ;
  wire  \inst_doa_mux_b3/B0_3 ;
  wire  \inst_doa_mux_b3/B1_0 ;
  wire  \inst_doa_mux_b3/B1_1 ;
  wire  \inst_doa_mux_b30/B0_0 ;
  wire  \inst_doa_mux_b30/B0_1 ;
  wire  \inst_doa_mux_b30/B0_2 ;
  wire  \inst_doa_mux_b30/B0_3 ;
  wire  \inst_doa_mux_b30/B1_0 ;
  wire  \inst_doa_mux_b30/B1_1 ;
  wire  \inst_doa_mux_b31/B0_0 ;
  wire  \inst_doa_mux_b31/B0_1 ;
  wire  \inst_doa_mux_b31/B0_2 ;
  wire  \inst_doa_mux_b31/B0_3 ;
  wire  \inst_doa_mux_b31/B1_0 ;
  wire  \inst_doa_mux_b31/B1_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b4/B0_2 ;
  wire  \inst_doa_mux_b4/B0_3 ;
  wire  \inst_doa_mux_b4/B1_0 ;
  wire  \inst_doa_mux_b4/B1_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b5/B0_2 ;
  wire  \inst_doa_mux_b5/B0_3 ;
  wire  \inst_doa_mux_b5/B1_0 ;
  wire  \inst_doa_mux_b5/B1_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b6/B0_2 ;
  wire  \inst_doa_mux_b6/B0_3 ;
  wire  \inst_doa_mux_b6/B1_0 ;
  wire  \inst_doa_mux_b6/B1_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b7/B0_2 ;
  wire  \inst_doa_mux_b7/B0_3 ;
  wire  \inst_doa_mux_b7/B1_0 ;
  wire  \inst_doa_mux_b7/B1_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b8/B0_2 ;
  wire  \inst_doa_mux_b8/B0_3 ;
  wire  \inst_doa_mux_b8/B1_0 ;
  wire  \inst_doa_mux_b8/B1_1 ;
  wire  \inst_doa_mux_b9/B0_0 ;
  wire  \inst_doa_mux_b9/B0_1 ;
  wire  \inst_doa_mux_b9/B0_2 ;
  wire  \inst_doa_mux_b9/B0_3 ;
  wire  \inst_doa_mux_b9/B1_0 ;
  wire  \inst_doa_mux_b9/B1_1 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i0_012;
  wire inst_doa_i0_013;
  wire inst_doa_i0_014;
  wire inst_doa_i0_015;
  wire inst_doa_i0_016;
  wire inst_doa_i0_017;
  wire inst_doa_i0_018;
  wire inst_doa_i0_019;
  wire inst_doa_i0_020;
  wire inst_doa_i0_021;
  wire inst_doa_i0_022;
  wire inst_doa_i0_023;
  wire inst_doa_i0_024;
  wire inst_doa_i0_025;
  wire inst_doa_i0_026;
  wire inst_doa_i0_027;
  wire inst_doa_i0_028;
  wire inst_doa_i0_029;
  wire inst_doa_i0_030;
  wire inst_doa_i0_031;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i1_009;
  wire inst_doa_i1_010;
  wire inst_doa_i1_011;
  wire inst_doa_i1_012;
  wire inst_doa_i1_013;
  wire inst_doa_i1_014;
  wire inst_doa_i1_015;
  wire inst_doa_i1_016;
  wire inst_doa_i1_017;
  wire inst_doa_i1_018;
  wire inst_doa_i1_019;
  wire inst_doa_i1_020;
  wire inst_doa_i1_021;
  wire inst_doa_i1_022;
  wire inst_doa_i1_023;
  wire inst_doa_i1_024;
  wire inst_doa_i1_025;
  wire inst_doa_i1_026;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i2_009;
  wire inst_doa_i2_010;
  wire inst_doa_i2_011;
  wire inst_doa_i2_012;
  wire inst_doa_i2_013;
  wire inst_doa_i2_014;
  wire inst_doa_i2_015;
  wire inst_doa_i2_016;
  wire inst_doa_i2_017;
  wire inst_doa_i2_018;
  wire inst_doa_i2_019;
  wire inst_doa_i2_020;
  wire inst_doa_i2_021;
  wire inst_doa_i2_022;
  wire inst_doa_i2_023;
  wire inst_doa_i2_024;
  wire inst_doa_i2_025;
  wire inst_doa_i2_026;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;
  wire inst_doa_i3_009;
  wire inst_doa_i3_010;
  wire inst_doa_i3_011;
  wire inst_doa_i3_012;
  wire inst_doa_i3_013;
  wire inst_doa_i3_014;
  wire inst_doa_i3_015;
  wire inst_doa_i3_016;
  wire inst_doa_i3_017;
  wire inst_doa_i3_018;
  wire inst_doa_i3_019;
  wire inst_doa_i3_020;
  wire inst_doa_i3_021;
  wire inst_doa_i3_022;
  wire inst_doa_i3_023;
  wire inst_doa_i3_024;
  wire inst_doa_i3_025;
  wire inst_doa_i3_026;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i4_003;
  wire inst_doa_i4_004;
  wire inst_doa_i4_005;
  wire inst_doa_i4_006;
  wire inst_doa_i4_007;
  wire inst_doa_i4_008;
  wire inst_doa_i5_000;
  wire inst_doa_i5_001;
  wire inst_doa_i5_002;
  wire inst_doa_i5_003;
  wire inst_doa_i5_004;
  wire inst_doa_i5_005;
  wire inst_doa_i5_006;
  wire inst_doa_i5_007;
  wire inst_doa_i5_008;
  wire inst_doa_i6_000;
  wire inst_doa_i6_001;
  wire inst_doa_i6_002;
  wire inst_doa_i6_003;
  wire inst_doa_i6_004;
  wire inst_doa_i6_005;
  wire inst_doa_i6_006;
  wire inst_doa_i6_007;
  wire inst_doa_i6_008;
  wire inst_doa_i7_000;
  wire inst_doa_i7_001;
  wire inst_doa_i7_002;
  wire inst_doa_i7_003;
  wire inst_doa_i7_004;
  wire inst_doa_i7_005;
  wire inst_doa_i7_006;
  wire inst_doa_i7_007;
  wire inst_doa_i7_008;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[10]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  reg_sr_as_w1 addra_pipe_b2 (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[2]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00000000000000000000000000000000000000000000000152633E03E6666666),
    .INITP_01(256'h000000000000000000000000000000000000000000B333333430049600000003),
    .INITP_02(256'h6666662B40D710143E9CC2928564B963C392894599321CA38000000000000000),
    .INITP_03(256'h49850162C00524CD5114004500155513FB00644CBA21641D0C30A55655A06F0E),
    .INIT_00(256'h3793139313931393139313931393139313931393139313931393139313931393),
    .INIT_01(256'h670B670B73EF13E32313831313179313E3231393971393736F0B232323231313),
    .INIT_02(256'h000000000000000000000000000000000000000000000000000000000000670B),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h2323232323232323232323232323232323232323232323232323238B238B0B13),
    .INIT_09(256'h83038303830B830B830B03038313172383131723630313170BEFEF8BEF138B23),
    .INIT_0A(256'h000000000000000B138B83038303830383038303830383038303830383038303),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h9402788484010000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h000000000000000000000000000000000000000000002CB4B40A30A4A4052094),
    .INIT_11(256'hB767000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h1383EF13931393B7B7EF13931393B7B7EFEF2313B737EF23136F1383EF231303),
    .INIT_13(256'h37936F2367638313376723B76FEF13EF13372323136FEF13EF13372323136F13),
    .INIT_14(256'h93EF1323231363936F131383E393232313933793B7EF231367131383EF231313),
    .INIT_15(256'h236303B39313B76393676F1333938303B393EF132323136393676F1383033333),
    .INIT_16(256'h83130383E31393E7138363836393B39393131313232323232337231367136723),
    .INIT_17(256'h0383038303830383038303830383038303830383038303838303036713038303),
    .INIT_18(256'h2313233723376303B76F9323672323232393B763139313371313136713830383),
    .INIT_19(256'h0383736383B76313236303B7EF132323136F136723B72313233723376303B767),
    .INIT_1A(256'h93231383376F13830323B7EF132323136703B76767138363EFEF231313376713),
    .INIT_1B(256'h133393B393EF139333133313EF932323239313636F1383EF238363239383EF23),
    .INIT_1C(256'h83038363931323B7372323136713671367136713671367138303833313EF1393),
    .INIT_1D(256'h23136F1383EF23136FE71383671383038363931323B7372323136FE713836713),
    .INIT_1E(256'h131383EFEFEFEFEFEFEFEFEF23136F13830313EF239313931393139313B73737),
    .INIT_1F(256'h1383EF67138303830383038363839393232323232323231367131383EF231367),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_008,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000038080000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000002210000000000),
    .INITP_02(256'h00000000012E0001B90C8101020FF000B4284420038760090000000000000000),
    .INITP_03(256'h200800080230028604C0063001800000700000299450408418E84AACAB77DA70),
    .INIT_00(256'h2007070707060606060505050504040404030303030202020201010101000000),
    .INIT_01(256'h40B240B2000002FC9782130303030202FE9782C20A0200000030939291908080),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000004062),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h969594939291909796959493929190979695949392919097969591A090205080),
    .INIT_09(256'h92929191915090509090925012020A5012020A108414020AE000006200009097),
    .INIT_0A(256'h000000000000000080A097979797969696969595959594949494939393939292),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0100000101000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000010100000101000001),
    .INIT_11(256'h0B40000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h02900002C203430A1B0002C203430A1B00F8D6820BC2009380008090F89380D2),
    .INIT_13(256'h1A82F89240CAA3820340D203F8080208021A939280F8080208021A9392800080),
    .INIT_14(256'h030082939280E50300800290CDC3D1D083C30BC30B0093804080029008938280),
    .INIT_15(256'hD0C5D2C3C38A0BE203400080FAE39092CB030082939280E603400080909232CA),
    .INIT_16(256'h928292904E0242C04212C413C6FB2B040202C58497929394950A9680400240D1),
    .INIT_17(256'h9796969696959595959494949493939393929292929191919091904080959494),
    .INIT_18(256'hD003910B920B8BD30BF8C3D04012101211C34308838302E3843B030080979797),
    .INIT_19(256'h929000C2D30B0D3AD780D30BF882939280F80240D70BD003910B920B8BD30B40),
    .INIT_1A(256'hC39380930BF8809092D30BF88293928040D20B4040809088F8089382801A4080),
    .INIT_1B(256'h8AC2CBC38B084202020A028A08829192930280A6088090089093CC90C3930893),
    .INIT_1C(256'h929290364202931A1A919280400240024002400240024080929290820A088202),
    .INIT_1D(256'h9280088090F89380F8C002134080929290364202931A1A919280F8C002134080),
    .INIT_1E(256'h800290080008F8080800F8F8938008809092020893C2030383030404021A0B0B),
    .INIT_1F(256'h8513F8408095959494929290CA130504929496979193958040800290F8938040),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_017,inst_doa_i0_016,inst_doa_i0_015,inst_doa_i0_014,inst_doa_i0_013,inst_doa_i0_012,inst_doa_i0_011,inst_doa_i0_010,inst_doa_i0_009}));
  // address_offset=0;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00000000000000000000000000000000000000000000000011A0D84200000000),
    .INITP_01(256'h0000000000000000000000000000000000000000013FFFC000066329FFFE0000),
    .INITP_02(256'hFFF80000080000100024020004A8810322090CC42A14E0CB0000000000000000),
    .INITP_03(256'h2000010211342208618030600C1004030100799E2411000800A0A80000400947),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h00810081047400A9BD11F11181004000A98111E1FF400004208000000000C000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'hF8F4F0ECE8E4E05C5854504C484440BCB8B4B0ACA8A4A01C1814040004008000),
    .INIT_09(256'h9080706050801080008100010101FF090151FF01820181FF0034F000C40080FC),
    .INIT_0A(256'h00000000000000000000F0E0D0C0B0A090807060504030201000F0E0D0C0B0A0),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0430A004E100B100001000F1008100009003A9810000B004C0504030B304C0E1),
    .INIT_13(256'h0001B73D0001FD0580002980C7640C6051000420C0C7F408F0E1000420C06040),
    .INIT_14(256'h04F0010420C0A97C8040FC30B5210139E1010001003004C000400030300461C0),
    .INIT_15(256'h2D010129010D00A97C00A04029FD3020210400010420C0A97C00A04030202921),
    .INIT_16(256'h500260704D21050101110101010526800001010104504C482400208000000031),
    .INIT_17(256'hC0B0A090807060504030201000F0E0D0C0B0A090807060501000010080203040),
    .INIT_18(256'h39042D002900010100671139003D41AD350100BDBD0101AB01F1110000F0E0D0),
    .INIT_19(256'h20300001010001098181F10093010420C0E3FC00B90039042D00290001010000),
    .INIT_1A(256'h0504C0310057403020210097010420C0003100000040300167000401C0000040),
    .INIT_1B(256'h09290D29059401A0290D2905F401242004A0C081644030103DF1013DFD01303D),
    .INIT_1C(256'h10203025C1B10400002420C0000000000000000000FC00401020302109049DA0),
    .INIT_1D(256'h20C0244030C704C077011101004010203025D1C10400002420C0770111010040),
    .INIT_1E(256'h400030C0B07457005474279704C0E44030200090044181000100085000000000),
    .INIT_1F(256'h012007008010203040506070CD20042050482004544C248000400030F704C000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_026,inst_doa_i0_025,inst_doa_i0_024,inst_doa_i0_023,inst_doa_i0_022,inst_doa_i0_021,inst_doa_i0_020,inst_doa_i0_019,inst_doa_i0_018}));
  // address_offset=0;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000045AADC0200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000008000000006634400000001),
    .INIT_02(256'h0000000008004010082402000428950922090CC40A54D08A0000000000000000),
    .INIT_03(256'h6005010A02643688458000600010040701086909304140D80800A2A4A947CB48),
    .INIT_04(256'h0800042001C248801044041000018001010684200020CB22A85A026400008012),
    .INIT_05(256'h40181008010002C1A088D08012080A008210002FE1205B080100501425B081B1),
    .INIT_06(256'h10003801128201242A900000C20D048C309A00649400000020060C0001005004),
    .INIT_07(256'h08010C0002102004805002010034001AC1C080404014000E0C0440000C000201),
    .INIT_08(256'h0022032560010495081D312442C0008D100101C012C2948C135C828008810004),
    .INIT_09(256'h080D0200A00001080B0040808140A91086040000131502088050100002200000),
    .INIT_0A(256'h0016480352080102421140000519028210284200088010080141282028800500),
    .INIT_0B(256'h00240000000000000000005641D4338302B080428100840120902040A1DB90AA),
    .INIT_0C(256'h0000000000000000000A843235A7001000649249249249249244887001D02108),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_027 (
    .addra(addra),
    .clka(clka),
    .dia({open_n195,open_n196,open_n197,open_n198,open_n199,open_n200,open_n201,1'b0,open_n202}),
    .rsta(rsta),
    .doa({open_n217,open_n218,open_n219,open_n220,open_n221,open_n222,open_n223,open_n224,inst_doa_i0_027}));
  // address_offset=0;data_offset=28;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000001A2CC0200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000002210000000001),
    .INIT_02(256'h0000000008000010002402000428C109220D0EC62244628B0000000000000000),
    .INIT_03(256'h4005010A1FB400C045800060001004030500690B3451408808A0AAA4A9478340),
    .INIT_04(256'h2800042001C24880104424100101800000008400002D5B468000007600048012),
    .INIT_05(256'h40181008010002C1A088D08012080A208210002FE000DB080100001421A091A1),
    .INIT_06(256'h00003805129201A022900000000D048C109A00649400000020060C0001005004),
    .INIT_07(256'h00000D000618A004800000001002101AC1000040401C100E0C0440000C000201),
    .INIT_08(256'h0032032561000095081D312442C10009101111A10EC7948C3B5E868000800004),
    .INIT_09(256'h00080B00A01401084300420481400900840804001B9580002050100003200004),
    .INIT_0A(256'h0016080352080102421140000519049010220200088010080141282029800100),
    .INIT_0B(256'h5A80000000000000000063011600C064C0F080428110944120902040A1DB9828),
    .INIT_0C(256'h000000000000000000307209C000020000000000000000000000618003466A0A),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_028 (
    .addra(addra),
    .clka(clka),
    .dia({open_n256,open_n257,open_n258,open_n259,open_n260,open_n261,open_n262,1'b0,open_n263}),
    .rsta(rsta),
    .doa({open_n278,open_n279,open_n280,open_n281,open_n282,open_n283,open_n284,open_n285,inst_doa_i0_028}));
  // address_offset=0;data_offset=29;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000005A2CC0200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000002212400000001),
    .INIT_02(256'h00000000080000100004222044A8050B22098C840000508A0000000000000000),
    .INIT_03(256'h4005010A0244260865800060001004070508610A241100980000A00000478A40),
    .INIT_04(256'h0800042001C24880104424100101802100008420002D5B4688530676400C8212),
    .INIT_05(256'h40181008010002C1A088D08012080A208210002FE000DB080100001401A001A0),
    .INIT_06(256'h000038000292018022904412000D048C109A00649400000020060C0001007004),
    .INIT_07(256'h00000C000218A004805000001022101AC1400040401C100F2E0440000C000201),
    .INIT_08(256'h00200325400044140110258162C1008D101111E10EC684CC335E848028914004),
    .INIT_09(256'h00080300A04400084B005A04C1408910860C04001B9582080050100003200004),
    .INIT_0A(256'h00040003520801021011400800104692100A4200080010080051088029800004),
    .INIT_0B(256'h7D100000000000000001E3533FD5F3EFDB853014C34094412090204001139028),
    .INIT_0C(256'h00000000000000000027FFFFF7FF020000000000000000000000FFF0035FFBFB),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_029 (
    .addra(addra),
    .clka(clka),
    .dia({open_n317,open_n318,open_n319,open_n320,open_n321,open_n322,open_n323,1'b0,open_n324}),
    .rsta(rsta),
    .doa({open_n339,open_n340,open_n341,open_n342,open_n343,open_n344,open_n345,open_n346,inst_doa_i0_029}));
  // address_offset=0;data_offset=30;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000005A8D80200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000002216800000001),
    .INIT_02(256'h00000000080000100004020004280103220C8E44020472CB0000000000000000),
    .INIT_03(256'h2000010A06D4160065800060001004040408290B3451409808A8EAA4A9478B40),
    .INIT_04(256'h2800062001E268C011462411010180000008842000204200A810007720048010),
    .INIT_05(256'h40191048812802C1A188D0C012080A208218243FE000DB084140001425A091A1),
    .INIT_06(256'h120138050292018022904000000D058C109A006494000002A0060C0001007024),
    .INIT_07(256'h08010D0006102004800001009022101AC08080504014000BA64440900C000001),
    .INIT_08(256'h00320320204144050105B1244080000800010180008310841A00828008810004),
    .INIT_09(256'h08080100A01001084B0048844140A110860400000B808000A040200002200000),
    .INIT_0A(256'h0016000352080102101160000519009010220200088010080011008009800400),
    .INIT_0B(256'h5E8400000000000000018C5337D5F6A55B8500940050BE4374912040A1DB90B8),
    .INIT_0C(256'h0000000000000000001FFBFFF6F8000000000000000000000000F7800097C348),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_030 (
    .addra(addra),
    .clka(clka),
    .dia({open_n378,open_n379,open_n380,open_n381,open_n382,open_n383,open_n384,1'b0,open_n385}),
    .rsta(rsta),
    .doa({open_n400,open_n401,open_n402,open_n403,open_n404,open_n405,open_n406,open_n407,inst_doa_i0_030}));
  // address_offset=0;data_offset=31;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000001A0D80200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000006630000000001),
    .INIT_02(256'h0000000008004010080402000428910322088C440A14608B0000000000000000),
    .INIT_03(256'h2000010A023406804580006000100400000020093451409808A8EAA4A947CB40),
    .INIT_04(256'h2800042001C2488010442410010180000000842000244B02A012027720000010),
    .INIT_05(256'h40181008010002C1A088D08012080A208210002FE000DB080100001425A091A1),
    .INIT_06(256'h100038050292018022904000000D048C109A00649400000020060C0001007004),
    .INIT_07(256'h08010D0006102004800000001022101AC1C08050401C100F2E4440800C000201),
    .INIT_08(256'h0032032021410485090D35A56080008C000111E1008314C41A00828008810004),
    .INIT_09(256'h08080900A05001084B00580441408910860C00000B8082082040000002210004),
    .INIT_0A(256'h0016C8035208010252114008051D4692102A420008801008011120A009800504),
    .INIT_0B(256'h0000000000000000000000000000000000D5805600D0944120902040A1DB98AA),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000004000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_031 (
    .addra(addra),
    .clka(clka),
    .dia({open_n439,open_n440,open_n441,open_n442,open_n443,open_n444,open_n445,1'b0,open_n446}),
    .rsta(rsta),
    .doa({open_n461,open_n462,open_n463,open_n464,open_n465,open_n466,open_n467,open_n468,inst_doa_i0_031}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h8B331110281128429142005100049198068121A8062AD2B4B49330C49312541C),
    .INITP_01(256'h20956A569ABEA8497925396AA8D34E0820668B4018DB60841517C568B1044145),
    .INITP_02(256'h88C7A822C8000800014A234800A37154528AF240010A666211131D4005588C03),
    .INITP_03(256'hB40C08B0195248252D63DF6FBB11C9ECE880C0410014400A00222C5756082424),
    .INIT_00(256'h13EF6F138303830383830313EFEF1363EF13E7136383EF232323231303830363),
    .INIT_01(256'h136713376F13830313EF239313931393139313B73713132337136FEF23136FEF),
    .INIT_02(256'h2323232323B7132323231367036F132393938383EF23136F132393938383EF23),
    .INIT_03(256'h23232323231393639393939333636393E313936F131363139363931393232323),
    .INIT_04(256'h13936393932393E393B3936393936FE3A3939383331303830383EF13931303EF),
    .INIT_05(256'h13631313236363333313136313E3B31323636F13136F936F1333131363636333),
    .INIT_06(256'h636F93339363639393E3331323636F33136F333313136313E3B31323636F93B3),
    .INIT_07(256'hB763EF231367133383038303830383038303831363E3B39323636F1323033313),
    .INIT_08(256'h1383133763EF23136F23E3EF6713038323B763EF132323136F03E3EF67138303),
    .INIT_09(256'h63B3133313B3939363339393B33313B313936763339363936393136F13E3EF67),
    .INIT_0A(256'h230323139303676313936393B36393136FA3936F23136F23932323236FB39313),
    .INIT_0B(256'h6F23133383336F93B313936F33B3B393136333931333B3B39313E33323032303),
    .INIT_0C(256'h9363136F9367E323933383336F2333330333676393939363B3636F2313B303B3),
    .INIT_0D(256'h9393039393636733E3631363139363131383938313136713E3B3138383B3B36F),
    .INIT_0E(256'h33636303836713E313639393B383B383B36F93631367E3136FA36763933363A3),
    .INIT_0F(256'h63EF932323232323131323136F9367336303936F93671363633383936F931367),
    .INIT_10(256'h2323232323132313671303830383038313E3EF931393136F1363333393EF1313),
    .INIT_11(256'h6363E38313139313236363136F139313931337B79313639313B3232323232323),
    .INIT_12(256'h6F13636F13E393831313636F1393131367130383038303830383038303833323),
    .INIT_13(256'h9393631313938363939303E393831393331333936F13136393136F13636F1363),
    .INIT_14(256'h636393039363139303939363E393039313B393B3936F1333E3939303E313936F),
    .INIT_15(256'h9313E39363936F136F93936F93138363936F13A3636313832393636393636393),
    .INIT_16(256'h139333639303E313E39313E39393E3936F03939313136393E39363936363936F),
    .INIT_17(256'h1323636F9363B3133313238363931333136393E3931323636F939363136F93EF),
    .INIT_18(256'h63936393E313931323636F1393631393636303039383EF23232313936313836F),
    .INIT_19(256'h13136F936F936F93136F1323636F1323636F932383B363336F9363B313333393),
    .INIT_1A(256'h83EF232323232323231323136F931393671383EF2323232323239323136FA36F),
    .INIT_1B(256'h13133767130383EF13EF23232323232313939313232323372313676F63676713),
    .INIT_1C(256'h1363B393B7671303B3639313B7636F13133783EF93139313133737EF1337EF23),
    .INIT_1D(256'hE39313673313638313931393676713033313671303B3931363B3B76713033313),
    .INIT_1E(256'h2323839303EFEF1313932393EF639383EF13EF13932323232323131323136713),
    .INIT_1F(256'h036713036F13032323232383930383EF13232323136F836F1303830383032323),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_008,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=1024;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h20000BE604226B385159FC114101D010050402000404C932000A1A33A0102861),
    .INITP_01(256'h400DDBE8E3FD13DFC5FF81F853ADCA3EB21BE4EFFD34FFFF5B879A9004809081),
    .INITP_02(256'h1A032825601202AC2AB14416C453FCA8311AF16DB72000003224230000002024),
    .INITP_03(256'h0861050046403000ED008CA651EA51762140001040091007EA4472B0EE098211),
    .INIT_00(256'h0208F88095959494929092020800828E0082C082C313081011D09104131312C5),
    .INIT_01(256'h8040820A08809092020893C2030383030404021A0B0282920B80F8F89380F8F8),
    .INIT_02(256'h90919295971CC4939496804022F88006FBC39023F89380F88006FBC39023F893),
    .INIT_03(256'h939495969702024B050285060328C03AC4063A00063C843DC4CAC4823A959697),
    .INIT_04(256'h3CC36A430280030D4E1E3ECC063A000847454222C58394939393080202859308),
    .INIT_05(256'h02810283003A4583028303AA83248203003AF82B3DF80600040203832A430883),
    .INIT_06(256'hBD00028383CD42420364438280BAF80203F883028303AA83248203003A000203),
    .INIT_07(256'h0B86F89380408082969695959595949492929003AA2403C3C0FAF88280230383),
    .INIT_08(256'h8090820A86F89380F894810840809290D40B87F882939280F8928208408090D2),
    .INIT_09(256'h338404C1C3833B3B7544038384B3CBB3CBFB40C9C383C5BBBC8303F882820840),
    .INIT_0A(256'h95D49483C3D440880383C0FBB3BD8303F8C7C3F81703F8D7C3D2D1D0F8C37B7B),
    .INIT_0B(256'hF81083C414C4F803C483C3F803C2C38B2B6404030303C2838B2B754497D496D4),
    .INIT_0C(256'h030B03F803400B80C383A3C3F88083C3A44340CAC30322BBC3FDF84083C364C3),
    .INIT_0D(256'h03C3E3C2830040C2CCCA433244C33243C4E3C2A3820340C2C7C38363E3C38300),
    .INIT_0E(256'hC2C3C2E3A340C24C83CBEBCB43E3C3E38300030B03404B43F8C740CAC3C38FC7),
    .INIT_0F(256'h80F8C49294959793C2829680F8C340C28BE383F8C34082B342C3E383F8C28240),
    .INIT_10(256'h9596979697C494804080959494929290028FF84202C28300026B020582F80284),
    .INIT_11(256'h3A83CF2382430202003AC3030005C40505021D8405A4FB428685949590919293),
    .INIT_12(256'hF834CBF834CB02234334C8000203030440809696969595959594949292900200),
    .INIT_13(256'h040372C24303630F0303633843638342838BC38B0003037103C3F834CBF834CB),
    .INIT_14(256'h72000363420EBB03620203EA788322C303C3CB43CBF83403AEC202D3CA030300),
    .INIT_15(256'h033408030003F802F80302F8C243D3CD03F80200BAC0026300033B0703700603),
    .INIT_16(256'h02C23BCA3AD38D0387C603090304060300D303C603348B030E03070375070300),
    .INIT_17(256'h8280BAF8C2238303030200D33BC383C303228324C302003A0003830E3CF842F8),
    .INIT_18(256'h6A43E30363838302003A0003830A3CC3EA2B93948393F891929342064AC6D6F8),
    .INIT_19(256'h2B0BF803F842F80334F802003AF88280BAF8C300E2423C03F882628303830203),
    .INIT_1A(256'h90F893979695949397839280F802C303408090F8939796959497839380F8C7F8),
    .INIT_1B(256'h82801A40809290F002F8939796959497020283839392910A968040F082404080),
    .INIT_1C(256'hAAC7BBC383408262438543BB1B80F880821A90F802030383821A1BF8821AF893),
    .INIT_1D(256'h89438340C28ACC5203030303404082A242AA4082E243BBAAC7BB834082A243BB),
    .INIT_1E(256'h1391900393F0F802030202F4004F83920084F805C49293949597C28296804002),
    .INIT_1F(256'hA240AA82F080921314905190031313F08282939280F852F08095949492921491),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_017,inst_doa_i1_016,inst_doa_i1_015,inst_doa_i1_014,inst_doa_i1_013,inst_doa_i1_012,inst_doa_i1_011,inst_doa_i1_010,inst_doa_i1_009}));
  // address_offset=1024;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h2A1FE42001C24884504420120100802101028408F9C4C22080400066200C0611),
    .INITP_01(256'h80181008010002C1A480508012080B600000002FE000D9000100401605A001B0),
    .INITP_02(256'h1000380503B501F714000407270D000D319A01649400400020260C0001007000),
    .INITP_03(256'h08010800040C00048000020100121008C980C0514014400F2E8400800C000001),
    .INIT_00(256'h02A027801020304050706002509402D5D40201020171502121393DB10111204D),
    .INIT_01(256'hC00001004040302001F00461210001001C8001000001012000C0F74704C017F7),
    .INIT_02(256'h585450240400014C48208000E0D740BCFDFD30E02704C07740BCFD0530E0C704),
    .INIT_03(256'h3034383C4001285D280080B43001810A81C0064080FA02425201820102E4E0DC),
    .INIT_04(256'h46013D0104B4C08117642201AC12B081AE060502520170605040F40128013064),
    .INIT_05(256'h010205FD6549033131FD000101AC31054149E7113DE70090803901FD38038235),
    .INIT_06(256'h49B08039010135FDFCB129052D49573901173131FD000101AC3105614930C035),
    .INIT_07(256'h00016704C0008039D0E0F000102030405060700001B43D052D49370531012580),
    .INIT_08(256'h40304100019704C097A181000040203021000177010420C0A7C1810000403041),
    .INIT_09(256'hC6300C35013D3DC1C13E3C01313D413D21FD00313101010D31010CA7C1813000),
    .INIT_0A(256'hC1D1C141410100B10001010D2D31013CD7AD0527B911D7B9413939398735310D),
    .INIT_0B(256'hE74611390239B73C310101373535350909C1390C003535351111413EC1F1C1E1),
    .INIT_0C(256'h003900D70000BD35053D013D87413931013D003DFD00FD353129374105390139),
    .INIT_0D(256'hFD05FD050101003901398141FD814101FDFD05FD056400010135050101393980),
    .INIT_0E(256'h3939010101000101050161613D01390139B0003900000101C7810031053101B9),
    .INIT_0F(256'h01F701504824044C01012080B7050029010101970500012D0129010187050500),
    .INIT_10(256'hA4A084605C01C8000080203040506070010107FD010202700049262901B70101),
    .INIT_11(256'h5D020101010501053D5DB9949022FE80AC030000FCFD2A0101496864D8D4D0CC),
    .INIT_12(256'h872259B742B905050112D540C08CB4000000405060708090A0B0C0D0E0F06101),
    .INIT_13(256'h24002941052405B5FCB801BD4101410535053909702400B92441270629578235),
    .INIT_14(256'h3135A40105B5EDA001010001B64101410529053D09B742388111090135FCA810),
    .INIT_15(256'h280AB590B58C37000700010711090135A8C7093D5D0105013D945DBD94B13560),
    .INIT_16(256'h01024D010A0131A03111B04540E0B5D4F0014011200635FCB5C035BCB1B5CC50),
    .INIT_17(256'h05315DE701342980390535015D1105390438FDBCFD05355D4080018242870353),
    .INIT_18(256'h0101B500BDFD0105315D508001824201293C201001304740383C030203110197),
    .INIT_19(256'h41418720F7FDC740024705315D2705315DF7052D013F5D3D3703BD2980393D00),
    .INIT_1A(256'h702730C4C0BCB8B404A0B00057FC0101000070C734C4C0BCB804B0B400F782E7),
    .INIT_1B(256'h41C00000006070F7E12734C4C0BCB804E1FC9001B4B0AC002000003701000000),
    .INIT_1C(256'h21013D01000005A1390181FD00015740B10030A70C040C013100002771005704),
    .INIT_1D(256'hB14105002911290110000000000065A129610045A13DFD41013D3F0025A139FD),
    .INIT_1E(256'h393D70311237130120024D02503D1212F001770101504C482404010120800000),
    .INIT_1F(256'h21007D214740203D3D353930314131D701010420C0870177802030405060253E),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_026,inst_doa_i1_025,inst_doa_i1_024,inst_doa_i1_023,inst_doa_i1_022,inst_doa_i1_021,inst_doa_i1_020,inst_doa_i1_019,inst_doa_i1_018}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0228230490AAAA05A490F95651AF850AA07B611274FC98B5F3114D5C46029205),
    .INITP_01(256'h640A622CAC2A0C0BA2706563015853A0B9601409921231554A560E00C03AC018),
    .INITP_02(256'h760A300264B54543A8168983002998E8161502802D011065624C03402A1BC21A),
    .INITP_03(256'hC1080000000000000000E7525C1458409F2B322CC861AA825503406035E4F355),
    .INIT_00(256'h8313EF63EF139313136F13EF639303EF03EF2393631313632323232323136713),
    .INIT_01(256'h33139313EF2313036723239323232313E3932323139323B76F03671383038303),
    .INIT_02(256'h6393139323832363130383B3931393EF03631383B7EF2323136F131323138303),
    .INIT_03(256'hB3038383232323238303B39313239393930383EF132323136FEF6F13830313EF),
    .INIT_04(256'h23136F13830323B39383836303B393138323232323938303EF132323136F1323),
    .INIT_05(256'hB76713836F13836F13836383EF2363239393938337EF23136F132393838337EF),
    .INIT_06(256'h13836F13838303EF13EF1363836393EF13EF132393EF1393EF23230323136703),
    .INIT_07(256'h23231323232393139323136F1383EF23232313232323131383036F2323932323),
    .INIT_08(256'h132323378303EF9333B79303830383EF93131323232323232313838303EF2323),
    .INIT_09(256'hEF13EF639313832323136703671313830383EF131393939323232323232323A3),
    .INIT_0A(256'h03931383EF23136FEF23239323231383EF6713130383EF1363836393EF132393),
    .INIT_0B(256'h13639313836FEF1367131383EFEF232323230333231313930323236303036313),
    .INIT_0C(256'h03EF2323232323136713671313830383EF13EF13EF239393139383EF13232323),
    .INIT_0D(256'h836F1383EF23136F6713130383038323639303EFEF13EF13EF13931393EF1313),
    .INIT_0E(256'h136713671313830383EF13EF13EF132323232393930383EF1323232313639313),
    .INIT_0F(256'h93939383EF132323232313231363936367131383EF6383EF23A3132333138323),
    .INIT_10(256'h232383231367136F6F23A3B3036713138303830383EF13EF23A3B31383EF1363),
    .INIT_11(256'h03830383038313EF638363EF139313136F13EF6303631383EF13EF6313232323),
    .INIT_12(256'h232393A393038383EF232323132323931393231367232323239303836F836713),
    .INIT_13(256'h23232313671313830383EF13EF13EF1393EF1323232313671383038323232323),
    .INIT_14(256'h23232323932393833763031393370313B7EF233383EFEFA3931383EF1393EF13),
    .INIT_15(256'h83EF13EF1393EF13232323136393836F93E3B3638383671313830383EFA39383),
    .INIT_16(256'hA393836F23836F23836F9383E393639367136363639367136713830383A39313),
    .INIT_17(256'h83138303038303838303630393931393B7EF3793EF232323232323232323136F),
    .INIT_18(256'h23239337670363139303B76FEF13E3A393139383EFE70383EF13E33313036F13),
    .INIT_19(256'h93B36FB363336713EF9367E3139333B36313E393136363936313931363636767),
    .INIT_1A(256'h13931393B7379313EF1337EF23232313136733EF33E3B36713EF6363936733EF),
    .INIT_1B(256'h610D6176726D76726FEF13EF13EF1393139313931393B73793EF13EF13931393),
    .INIT_1C(256'h0021726F20726E656155327431740D6F33636F6820752E6920610D0D742E6920),
    .INIT_1D(256'h0204020302050203020402030200006338343000433834306574006D002E6473),
    .INIT_1E(256'h0204020302050203020402030207020302040203020502030204020302060203),
    .INIT_1F(256'h65536965646820202D007C0A4C28020302040203020502030204020302060203),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_008,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  // address_offset=2048;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0092502221510481092DF4B5219E1884856B10E1903954400820FA8008010800),
    .INITP_01(256'h0C000D08005061064900980440008B10670FFBFF898882883800100013E16004),
    .INITP_02(256'h4000480157201002520DF40A573B5692002A400008804188019420B001900504),
    .INITP_03(256'hE8A000000000000000006306101449468DD483520CB05145229C3A80E6DECCC2),
    .INIT_00(256'h9002008AF802C203820002008C8294F892009384B302038597909192938040BA),
    .INIT_01(256'h828A0382F89380124012D10311100703CDC3D0D1C303CD0BF894408094949292),
    .INIT_02(256'hCFC282FB07231081C312D2C34B0383F812CB82CB0BF0939280F0808210839092),
    .INIT_03(256'hF392131315D1169090D3C3038B05F3FB032323F082939280F8F0F080909202F0),
    .INIT_04(256'h9380F080909211FBE313138ED3C3CB032316159051031313F082939280F08011),
    .INIT_05(256'h0B408090F08090F88090C713F08D208DEBCBC3AB0BF09380F0808DC390AB0BF0),
    .INIT_06(256'h0313F880929092F042F802CA138C03F80200020503F80282F0919312928040EA),
    .INIT_07(256'h97938294929302C3029180F88090F89596508311949303809393F81615035112),
    .INIT_08(256'h020517139494F0430313C312121313F80282C313111015161203939393F89596),
    .INIT_09(256'h0002F8C2FB82A393928040124080029292900003030302031514051410171605),
    .INIT_0A(256'hE3830313F09380F8F016150351120313F04080029290F802C8138A03F8020503),
    .INIT_0B(256'h80C8FB03A3F8F04240800290F8F0D591D6109383D6030BC3E3901104D3D38FBB),
    .INIT_0C(256'h12F09394959697804002408002929290F0420002F805F3FB028223F082919293),
    .INIT_0D(256'hA3F88090F09380F840800294929290148A0313F8F08200420042028302F80284),
    .INIT_0E(256'h804002408002929290F802F04200021516905182031313F08291929380CBFB03),
    .INIT_0F(256'h7A840322F00497939495829680CF03C040800290F8C213F8858503968B03A393),
    .INIT_10(256'h97921395804002F8F81605CBA34080029494929290F0C2F816054A02A3F8024B),
    .INIT_11(256'h95949492929002F8C2138DF0020203C20002F80512CE8494F802F8C285939496),
    .INIT_12(256'h10170302FB939393F891929382979602C30295804095969051839393F8D44080),
    .INIT_13(256'h91929380408002929290F802F042F80282F08291929380408092929015161112),
    .INIT_14(256'h16D01591031643130B0CD323C30394C30BF012C213F0F002FB4223F80282F082),
    .INIT_15(256'h23F042F80282F08291929380C5FBA3F8833943431293408002929290F002F323),
    .INIT_16(256'h82FBA3F89113F8109300F3A3CB03C4034002C5E4C4034002408092929002FB02),
    .INIT_17(256'h954295959594949290920D920562858502F00C84F096929394959790919380F8),
    .INIT_18(256'h97D1830B40928202C3D30BF8F8028B05FBFB8423F0C01213F80271C20512F080),
    .INIT_19(256'h4102F802EC0240C2F841404B2B6BB2C2F302354B0B2C3D03060282C3E3A04040),
    .INIT_1A(256'h030304041A0B0202F8821AE891929302804002F802AC0240C2F8A6E5414002F8),
    .INIT_1B(256'hB90536AFB4322FB4F8F802F842F842C20303030304041A0B02F842F842C20303),
    .INIT_1C(256'h0090B9B1123ABA3237A700B000B0053919371032063A17B7B9B905059097B7B9),
    .INIT_1D(256'h808080808080808080808080808000B29C1A1800A29C1A18003400B00017B7B4),
    .INIT_1E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1F(256'h36BCB7B990B910161000901014A7808080808080808080808080808080808080),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_017,inst_doa_i2_016,inst_doa_i2_015,inst_doa_i2_014,inst_doa_i2_013,inst_doa_i2_012,inst_doa_i2_011,inst_doa_i2_010,inst_doa_i2_009}));
  // address_offset=2048;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00320320014864040808210060800008000101C0188240C41A02880008904805),
    .INITP_01(256'h08080900A056000C4A00520C01401900C60C00120B808048404020C880210000),
    .INITP_02(256'h00044002520801024218000000504080102A4200080010000111202008800001),
    .INITP_03(256'h528400000000000000014A533481D3A740A124D4101094400010204C010190A8),
    .INIT_00(256'hB001B08103010220D28000402611114730002C012D0030814CC8A4A0844000FD),
    .INIT_01(256'h3D0DF0FD7704C010003C3D200000B81CB9213D3D01F00100C70200C0708090A0),
    .INIT_02(256'h012171FDB4E038B9B10001390DF0FD271001015100370420C0F7402138B13001),
    .INIT_03(256'h3520E1103D353935301139F00DBD05C151D5D117010420C0A717A74030200117),
    .INIT_04(256'h04C0274030203C35FD10E13D01390DF0D53D3D353951516167010420C0D7403C),
    .INIT_05(256'h00004030474030F740300100C701BC3D4141FD51003704C087403D05305100D7),
    .INIT_06(256'h5120A7401030207701570181C1BD04C701B011BD109701016724040020C00051),
    .INIT_07(256'h34440140A084040101A440374030773939315135B904F8C06151273D35203938),
    .INIT_08(256'h11C129003040C3213D00F18191A1B1538C0101BDB5A53131B951705060073C38),
    .INIT_09(256'hA01167013D01D10420C0000000C00090A0B0F061000001018181818145C581C1),
    .INIT_0A(256'hD10104002304C027833D352039385120E30040002030270181C1BD049701BD10),
    .INIT_0B(256'hC0B93D04D1A763010040003047D339353135113135F00D51D53139396151313D),
    .INIT_0C(256'h00F328482420048000FC0040001020300301401187BD09C10101D19301242004),
    .INIT_0D(256'hD1A740301304C00700800040506070813DF8C1B7430230013001003011970101),
    .INIT_0E(256'hC000FC0040001020302701B301F0113D3D3539015161515301242004C0B93D08),
    .INIT_0F(256'h3D0104D12301044C48240120803D088100400030C7010077B9B508B93504D904),
    .INIT_10(256'h045000248000007727BDB939020080003040506070530207A5BD3D010217013D),
    .INIT_11(256'h203040506070010701008177010220D2A000B781004A1111D3049701014C4820),
    .INIT_12(256'hB525513DF9203010B33C38340104202801012480003D3D353951615177020080),
    .INIT_13(256'h242004C00040001020306301C301370101F301242004C000805060703D3DB981),
    .INIT_14(256'h3D35393551350561003E01F97100117100F3A9299133633DF90125070101C301),
    .INIT_15(256'h2513018701014301242004C00105255701B52D2DA151004000102030C33D0525),
    .INIT_16(256'h3DF52527BD01573D91900925BD0CBD080000812DBD0400FC00401020303DF900),
    .INIT_17(256'h5002304060708090B0A0D9720CF9720100F300012350A05C58544CC8A48440E7),
    .INIT_18(256'h3D3D710000513DFC7171000797025DBDF90D01D523013121D702292AB151E3C0),
    .INIT_19(256'h002C772C01280001D7000081050535313100AD0505302D0481FC010181810000),
    .INIT_1A(256'h4000109000000140F3C1003724200400C0002C8728812C0001E7010100002847),
    .INIT_1B(256'h5A081BD9DC1C5DDCE727D0B701330141B100E10010900000E197011301212100),
    .INIT_1C(256'h00881958191C9948190B00DC00DC001BC89C5C1B0288C8999D9A0800105B999D),
    .INIT_1D(256'h0000000000000000000000000000009998CDCC009190CDCC0019009A008B9D1D),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h021C19181359080814008B170015000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_026,inst_doa_i2_025,inst_doa_i2_024,inst_doa_i2_023,inst_doa_i2_022,inst_doa_i2_021,inst_doa_i2_020,inst_doa_i2_019,inst_doa_i2_018}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00000000000000000000A595E7FA000A0036DB6DB6DB6DB6DB647B244158418B),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0265384840002E5520470A74652D796879203236200A64622E6420202030314A),
    .INIT_01(256'h0101040101040101040101C42C00017600696963672F2D692E2F2E000001FB00),
    .INIT_02(256'h0204010104010104010104010104010204010104010104010204010104010104),
    .INIT_03(256'h0000000001320001040401010401020401020401010401010401040401010401),
    .INIT_04(256'h696E652F767672662F626376722F2E2E0000B4880002021C0000250311110000),
    .INIT_05(256'h00000000000000000031205563696C776E336965736C2D2D756C2F76696C2D2D),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_008,inst_doa_i3_007,inst_doa_i3_006,inst_doa_i3_005,inst_doa_i3_004,inst_doa_i3_003,inst_doa_i3_002,inst_doa_i3_001,inst_doa_i3_000}));
  // address_offset=3072;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000002EB553FBDF1039C00002002000082080057BE0BAC24001),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000007070700191494A100B2303A103AB9A19890190090BA1297102E17191B3A),
    .INIT_01(256'h0104808104808104800104800102009700B9B337B1B6B3B99717178000808780),
    .INIT_02(256'h0480010480810480810480810480810480810480010480810480010480810480),
    .INIT_03(256'h38209E443C010111008081048081048081048081048001048081048081048081),
    .INIT_04(256'hB9B317B49717B4B4B1B31796B417179700000016000080000000878700000067),
    .INIT_05(256'h00000000000000000097199080B1B3B73599B999BA34B7B334B2B119B731BA33),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_017,inst_doa_i3_016,inst_doa_i3_015,inst_doa_i3_014,inst_doa_i3_013,inst_doa_i3_012,inst_doa_i3_011,inst_doa_i3_010,inst_doa_i3_009}));
  // address_offset=3072;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000BEE83B187003406000000000000000000597000928168),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h1100000000000B0891900058199A1C88DA1B4C0B0C00C91A19094808080C881B),
    .INIT_01(256'h4001C04001C04001C04101C0C000001459988B9BD89AD8988BCB8B8040400340),
    .INIT_02(256'h01C04001C04001C04101C04001C04101C04001C04001C04001C04001C04001C0),
    .INIT_03(256'h8C8C8B8B8C00C00040404001C04001C04001C04001C04001C04001C04001C040),
    .INIT_04(256'h988BDC5B1459DCD99BD85BD9DCCB8B8B0000000000017800000044864484608C),
    .INIT_05(256'h0000000000000000000CCBD091D90B4BDB4B988BD858D9D81B8B5D4C8B5ADB5B),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_026,inst_doa_i3_025,inst_doa_i3_024,inst_doa_i3_023,inst_doa_i3_022,inst_doa_i3_021,inst_doa_i3_020,inst_doa_i3_019,inst_doa_i3_018}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i4_008,inst_doa_i4_007,inst_doa_i4_006,inst_doa_i4_005,inst_doa_i4_004,inst_doa_i4_003,inst_doa_i4_002,inst_doa_i4_001,inst_doa_i4_000}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i5_008,inst_doa_i5_007,inst_doa_i5_006,inst_doa_i5_005,inst_doa_i5_004,inst_doa_i5_003,inst_doa_i5_002,inst_doa_i5_001,inst_doa_i5_000}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i6_008,inst_doa_i6_007,inst_doa_i6_006,inst_doa_i6_005,inst_doa_i6_004,inst_doa_i6_003,inst_doa_i6_002,inst_doa_i6_001,inst_doa_i6_000}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i7_008,inst_doa_i7_007,inst_doa_i7_006,inst_doa_i7_005,inst_doa_i7_004,inst_doa_i7_003,inst_doa_i7_002,inst_doa_i7_001,inst_doa_i7_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b0/B0_2 ),
    .i1(\inst_doa_mux_b0/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b1/B0_2 ),
    .i1(\inst_doa_mux_b1/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i1_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_1  (
    .i0(inst_doa_i2_010),
    .i1(inst_doa_i3_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_2 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_3 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b10/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b10/B0_2 ),
    .i1(\inst_doa_mux_b10/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b10/B1_0 ),
    .i1(\inst_doa_mux_b10/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i1_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_1  (
    .i0(inst_doa_i2_011),
    .i1(inst_doa_i3_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_2 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_3 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b11/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b11/B0_2 ),
    .i1(\inst_doa_mux_b11/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b11/B1_0 ),
    .i1(\inst_doa_mux_b11/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_0  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i1_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_1  (
    .i0(inst_doa_i2_012),
    .i1(inst_doa_i3_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i5_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_2 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_3 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b12/B0_0 ),
    .i1(\inst_doa_mux_b12/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b12/B0_2 ),
    .i1(\inst_doa_mux_b12/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b12/B1_0 ),
    .i1(\inst_doa_mux_b12/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[12]));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_0  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i1_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_1  (
    .i0(inst_doa_i2_013),
    .i1(inst_doa_i3_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i5_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_2 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_3 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b13/B0_0 ),
    .i1(\inst_doa_mux_b13/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b13/B0_2 ),
    .i1(\inst_doa_mux_b13/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b13/B1_0 ),
    .i1(\inst_doa_mux_b13/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[13]));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_0  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i1_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_1  (
    .i0(inst_doa_i2_014),
    .i1(inst_doa_i3_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i5_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_2 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_3 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b14/B0_0 ),
    .i1(\inst_doa_mux_b14/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b14/B0_2 ),
    .i1(\inst_doa_mux_b14/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b14/B1_0 ),
    .i1(\inst_doa_mux_b14/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[14]));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_0  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i1_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_1  (
    .i0(inst_doa_i2_015),
    .i1(inst_doa_i3_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i5_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_2 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_3 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b15/B0_0 ),
    .i1(\inst_doa_mux_b15/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b15/B0_2 ),
    .i1(\inst_doa_mux_b15/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b15/B1_0 ),
    .i1(\inst_doa_mux_b15/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[15]));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_0  (
    .i0(inst_doa_i0_016),
    .i1(inst_doa_i1_016),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_0 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_1  (
    .i0(inst_doa_i2_016),
    .i1(inst_doa_i3_016),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_1 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i5_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_2 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_3 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b16/B0_0 ),
    .i1(\inst_doa_mux_b16/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b16/B1_0 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b16/B0_2 ),
    .i1(\inst_doa_mux_b16/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b16/B1_1 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b16/B1_0 ),
    .i1(\inst_doa_mux_b16/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[16]));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_0  (
    .i0(inst_doa_i0_017),
    .i1(inst_doa_i1_017),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_0 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_1  (
    .i0(inst_doa_i2_017),
    .i1(inst_doa_i3_017),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_1 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i5_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_2 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_3 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b17/B0_0 ),
    .i1(\inst_doa_mux_b17/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b17/B1_0 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b17/B0_2 ),
    .i1(\inst_doa_mux_b17/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b17/B1_1 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b17/B1_0 ),
    .i1(\inst_doa_mux_b17/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[17]));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_0  (
    .i0(inst_doa_i0_018),
    .i1(inst_doa_i1_018),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_0 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_1  (
    .i0(inst_doa_i2_018),
    .i1(inst_doa_i3_018),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_1 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_2 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_3 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b18/B0_0 ),
    .i1(\inst_doa_mux_b18/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b18/B1_0 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b18/B0_2 ),
    .i1(\inst_doa_mux_b18/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b18/B1_1 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b18/B1_0 ),
    .i1(\inst_doa_mux_b18/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[18]));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_0  (
    .i0(inst_doa_i0_019),
    .i1(inst_doa_i1_019),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_0 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_1  (
    .i0(inst_doa_i2_019),
    .i1(inst_doa_i3_019),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_1 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_2 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_3 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b19/B0_0 ),
    .i1(\inst_doa_mux_b19/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b19/B1_0 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b19/B0_2 ),
    .i1(\inst_doa_mux_b19/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b19/B1_1 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b19/B1_0 ),
    .i1(\inst_doa_mux_b19/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[19]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b2/B0_2 ),
    .i1(\inst_doa_mux_b2/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(\inst_doa_mux_b2/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_0  (
    .i0(inst_doa_i0_020),
    .i1(inst_doa_i1_020),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_0 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_1  (
    .i0(inst_doa_i2_020),
    .i1(inst_doa_i3_020),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_1 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_2 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_3 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b20/B0_0 ),
    .i1(\inst_doa_mux_b20/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b20/B1_0 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b20/B0_2 ),
    .i1(\inst_doa_mux_b20/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b20/B1_1 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b20/B1_0 ),
    .i1(\inst_doa_mux_b20/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[20]));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_0  (
    .i0(inst_doa_i0_021),
    .i1(inst_doa_i1_021),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_0 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_1  (
    .i0(inst_doa_i2_021),
    .i1(inst_doa_i3_021),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_1 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i5_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_2 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_3 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b21/B0_0 ),
    .i1(\inst_doa_mux_b21/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b21/B1_0 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b21/B0_2 ),
    .i1(\inst_doa_mux_b21/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b21/B1_1 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b21/B1_0 ),
    .i1(\inst_doa_mux_b21/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[21]));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_0  (
    .i0(inst_doa_i0_022),
    .i1(inst_doa_i1_022),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_0 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_1  (
    .i0(inst_doa_i2_022),
    .i1(inst_doa_i3_022),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_1 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i5_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_2 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_3 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b22/B0_0 ),
    .i1(\inst_doa_mux_b22/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b22/B1_0 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b22/B0_2 ),
    .i1(\inst_doa_mux_b22/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b22/B1_1 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b22/B1_0 ),
    .i1(\inst_doa_mux_b22/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[22]));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_0  (
    .i0(inst_doa_i0_023),
    .i1(inst_doa_i1_023),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_0 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_1  (
    .i0(inst_doa_i2_023),
    .i1(inst_doa_i3_023),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_1 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i5_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_2 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_3 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b23/B0_0 ),
    .i1(\inst_doa_mux_b23/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b23/B1_0 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b23/B0_2 ),
    .i1(\inst_doa_mux_b23/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b23/B1_1 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b23/B1_0 ),
    .i1(\inst_doa_mux_b23/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[23]));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_0  (
    .i0(inst_doa_i0_024),
    .i1(inst_doa_i1_024),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_0 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_1  (
    .i0(inst_doa_i2_024),
    .i1(inst_doa_i3_024),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_1 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i5_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_2 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_3 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b24/B0_0 ),
    .i1(\inst_doa_mux_b24/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b24/B1_0 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b24/B0_2 ),
    .i1(\inst_doa_mux_b24/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b24/B1_1 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b24/B1_0 ),
    .i1(\inst_doa_mux_b24/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[24]));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_0  (
    .i0(inst_doa_i0_025),
    .i1(inst_doa_i1_025),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_0 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_1  (
    .i0(inst_doa_i2_025),
    .i1(inst_doa_i3_025),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_1 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i5_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_2 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_3 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b25/B0_0 ),
    .i1(\inst_doa_mux_b25/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b25/B1_0 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b25/B0_2 ),
    .i1(\inst_doa_mux_b25/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b25/B1_1 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b25/B1_0 ),
    .i1(\inst_doa_mux_b25/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[25]));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_0  (
    .i0(inst_doa_i0_026),
    .i1(inst_doa_i1_026),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_0 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_1  (
    .i0(inst_doa_i2_026),
    .i1(inst_doa_i3_026),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_1 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i5_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_2 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_3 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b26/B0_0 ),
    .i1(\inst_doa_mux_b26/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b26/B1_0 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b26/B0_2 ),
    .i1(\inst_doa_mux_b26/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b26/B1_1 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b26/B1_0 ),
    .i1(\inst_doa_mux_b26/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[26]));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_0  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_0 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_1  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_1 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_2  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_2 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_3  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_3 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b27/B0_0 ),
    .i1(\inst_doa_mux_b27/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b27/B1_0 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b27/B0_2 ),
    .i1(\inst_doa_mux_b27/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b27/B1_1 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b27/B1_0 ),
    .i1(\inst_doa_mux_b27/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[27]));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_0  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_0 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_1  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_1 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_2  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_2 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_3  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_3 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b28/B0_0 ),
    .i1(\inst_doa_mux_b28/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b28/B1_0 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b28/B0_2 ),
    .i1(\inst_doa_mux_b28/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b28/B1_1 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b28/B1_0 ),
    .i1(\inst_doa_mux_b28/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[28]));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_0  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_0 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_1  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_1 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_2  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_2 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_3  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_3 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b29/B0_0 ),
    .i1(\inst_doa_mux_b29/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b29/B1_0 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b29/B0_2 ),
    .i1(\inst_doa_mux_b29/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b29/B1_1 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b29/B1_0 ),
    .i1(\inst_doa_mux_b29/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[29]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i5_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b3/B0_2 ),
    .i1(\inst_doa_mux_b3/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b3/B1_0 ),
    .i1(\inst_doa_mux_b3/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_0  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_0 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_1  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_1 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_2  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_2 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_3  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_3 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b30/B0_0 ),
    .i1(\inst_doa_mux_b30/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b30/B1_0 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b30/B0_2 ),
    .i1(\inst_doa_mux_b30/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b30/B1_1 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b30/B1_0 ),
    .i1(\inst_doa_mux_b30/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[30]));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_0  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_0 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_1  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_1 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_2  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_2 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_3  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_3 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b31/B0_0 ),
    .i1(\inst_doa_mux_b31/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b31/B1_0 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b31/B0_2 ),
    .i1(\inst_doa_mux_b31/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b31/B1_1 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b31/B1_0 ),
    .i1(\inst_doa_mux_b31/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[31]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i5_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b4/B0_2 ),
    .i1(\inst_doa_mux_b4/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b4/B1_0 ),
    .i1(\inst_doa_mux_b4/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i5_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b5/B0_2 ),
    .i1(\inst_doa_mux_b5/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b5/B1_0 ),
    .i1(\inst_doa_mux_b5/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i5_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b6/B0_2 ),
    .i1(\inst_doa_mux_b6/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b6/B1_0 ),
    .i1(\inst_doa_mux_b6/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i5_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b7/B0_2 ),
    .i1(\inst_doa_mux_b7/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b7/B1_0 ),
    .i1(\inst_doa_mux_b7/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i5_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b8/B0_2 ),
    .i1(\inst_doa_mux_b8/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b8/B1_0 ),
    .i1(\inst_doa_mux_b8/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i1_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_1  (
    .i0(inst_doa_i2_009),
    .i1(inst_doa_i3_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_2 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_3 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b9/B0_0 ),
    .i1(\inst_doa_mux_b9/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b9/B0_2 ),
    .i1(\inst_doa_mux_b9/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b9/B1_0 ),
    .i1(\inst_doa_mux_b9/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[9]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

