// Verilog netlist created by TD v4.3.633
// Sat Aug  1 16:33:21 2020

`timescale 1ns / 1ps
module rom  // al_ip/rom.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [12:0] addra;  // al_ip/rom.v(18)
  input clka;  // al_ip/rom.v(19)
  input rsta;  // al_ip/rom.v(20)
  output [31:0] doa;  // al_ip/rom.v(16)

  wire [0:2] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B0_2 ;
  wire  \inst_doa_mux_b0/B0_3 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b0/B1_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B0_2 ;
  wire  \inst_doa_mux_b1/B0_3 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b1/B1_1 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B0_1 ;
  wire  \inst_doa_mux_b10/B0_2 ;
  wire  \inst_doa_mux_b10/B0_3 ;
  wire  \inst_doa_mux_b10/B1_0 ;
  wire  \inst_doa_mux_b10/B1_1 ;
  wire  \inst_doa_mux_b11/B0_0 ;
  wire  \inst_doa_mux_b11/B0_1 ;
  wire  \inst_doa_mux_b11/B0_2 ;
  wire  \inst_doa_mux_b11/B0_3 ;
  wire  \inst_doa_mux_b11/B1_0 ;
  wire  \inst_doa_mux_b11/B1_1 ;
  wire  \inst_doa_mux_b12/B0_0 ;
  wire  \inst_doa_mux_b12/B0_1 ;
  wire  \inst_doa_mux_b12/B0_2 ;
  wire  \inst_doa_mux_b12/B0_3 ;
  wire  \inst_doa_mux_b12/B1_0 ;
  wire  \inst_doa_mux_b12/B1_1 ;
  wire  \inst_doa_mux_b13/B0_0 ;
  wire  \inst_doa_mux_b13/B0_1 ;
  wire  \inst_doa_mux_b13/B0_2 ;
  wire  \inst_doa_mux_b13/B0_3 ;
  wire  \inst_doa_mux_b13/B1_0 ;
  wire  \inst_doa_mux_b13/B1_1 ;
  wire  \inst_doa_mux_b14/B0_0 ;
  wire  \inst_doa_mux_b14/B0_1 ;
  wire  \inst_doa_mux_b14/B0_2 ;
  wire  \inst_doa_mux_b14/B0_3 ;
  wire  \inst_doa_mux_b14/B1_0 ;
  wire  \inst_doa_mux_b14/B1_1 ;
  wire  \inst_doa_mux_b15/B0_0 ;
  wire  \inst_doa_mux_b15/B0_1 ;
  wire  \inst_doa_mux_b15/B0_2 ;
  wire  \inst_doa_mux_b15/B0_3 ;
  wire  \inst_doa_mux_b15/B1_0 ;
  wire  \inst_doa_mux_b15/B1_1 ;
  wire  \inst_doa_mux_b16/B0_0 ;
  wire  \inst_doa_mux_b16/B0_1 ;
  wire  \inst_doa_mux_b16/B0_2 ;
  wire  \inst_doa_mux_b16/B0_3 ;
  wire  \inst_doa_mux_b16/B1_0 ;
  wire  \inst_doa_mux_b16/B1_1 ;
  wire  \inst_doa_mux_b17/B0_0 ;
  wire  \inst_doa_mux_b17/B0_1 ;
  wire  \inst_doa_mux_b17/B0_2 ;
  wire  \inst_doa_mux_b17/B0_3 ;
  wire  \inst_doa_mux_b17/B1_0 ;
  wire  \inst_doa_mux_b17/B1_1 ;
  wire  \inst_doa_mux_b18/B0_0 ;
  wire  \inst_doa_mux_b18/B0_1 ;
  wire  \inst_doa_mux_b18/B0_2 ;
  wire  \inst_doa_mux_b18/B0_3 ;
  wire  \inst_doa_mux_b18/B1_0 ;
  wire  \inst_doa_mux_b18/B1_1 ;
  wire  \inst_doa_mux_b19/B0_0 ;
  wire  \inst_doa_mux_b19/B0_1 ;
  wire  \inst_doa_mux_b19/B0_2 ;
  wire  \inst_doa_mux_b19/B0_3 ;
  wire  \inst_doa_mux_b19/B1_0 ;
  wire  \inst_doa_mux_b19/B1_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b2/B0_2 ;
  wire  \inst_doa_mux_b2/B0_3 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b2/B1_1 ;
  wire  \inst_doa_mux_b20/B0_0 ;
  wire  \inst_doa_mux_b20/B0_1 ;
  wire  \inst_doa_mux_b20/B0_2 ;
  wire  \inst_doa_mux_b20/B0_3 ;
  wire  \inst_doa_mux_b20/B1_0 ;
  wire  \inst_doa_mux_b20/B1_1 ;
  wire  \inst_doa_mux_b21/B0_0 ;
  wire  \inst_doa_mux_b21/B0_1 ;
  wire  \inst_doa_mux_b21/B0_2 ;
  wire  \inst_doa_mux_b21/B0_3 ;
  wire  \inst_doa_mux_b21/B1_0 ;
  wire  \inst_doa_mux_b21/B1_1 ;
  wire  \inst_doa_mux_b22/B0_0 ;
  wire  \inst_doa_mux_b22/B0_1 ;
  wire  \inst_doa_mux_b22/B0_2 ;
  wire  \inst_doa_mux_b22/B0_3 ;
  wire  \inst_doa_mux_b22/B1_0 ;
  wire  \inst_doa_mux_b22/B1_1 ;
  wire  \inst_doa_mux_b23/B0_0 ;
  wire  \inst_doa_mux_b23/B0_1 ;
  wire  \inst_doa_mux_b23/B0_2 ;
  wire  \inst_doa_mux_b23/B0_3 ;
  wire  \inst_doa_mux_b23/B1_0 ;
  wire  \inst_doa_mux_b23/B1_1 ;
  wire  \inst_doa_mux_b24/B0_0 ;
  wire  \inst_doa_mux_b24/B0_1 ;
  wire  \inst_doa_mux_b24/B0_2 ;
  wire  \inst_doa_mux_b24/B0_3 ;
  wire  \inst_doa_mux_b24/B1_0 ;
  wire  \inst_doa_mux_b24/B1_1 ;
  wire  \inst_doa_mux_b25/B0_0 ;
  wire  \inst_doa_mux_b25/B0_1 ;
  wire  \inst_doa_mux_b25/B0_2 ;
  wire  \inst_doa_mux_b25/B0_3 ;
  wire  \inst_doa_mux_b25/B1_0 ;
  wire  \inst_doa_mux_b25/B1_1 ;
  wire  \inst_doa_mux_b26/B0_0 ;
  wire  \inst_doa_mux_b26/B0_1 ;
  wire  \inst_doa_mux_b26/B0_2 ;
  wire  \inst_doa_mux_b26/B0_3 ;
  wire  \inst_doa_mux_b26/B1_0 ;
  wire  \inst_doa_mux_b26/B1_1 ;
  wire  \inst_doa_mux_b27/B0_0 ;
  wire  \inst_doa_mux_b27/B0_1 ;
  wire  \inst_doa_mux_b27/B0_2 ;
  wire  \inst_doa_mux_b27/B0_3 ;
  wire  \inst_doa_mux_b27/B1_0 ;
  wire  \inst_doa_mux_b27/B1_1 ;
  wire  \inst_doa_mux_b28/B0_0 ;
  wire  \inst_doa_mux_b28/B0_1 ;
  wire  \inst_doa_mux_b28/B0_2 ;
  wire  \inst_doa_mux_b28/B0_3 ;
  wire  \inst_doa_mux_b28/B1_0 ;
  wire  \inst_doa_mux_b28/B1_1 ;
  wire  \inst_doa_mux_b29/B0_0 ;
  wire  \inst_doa_mux_b29/B0_1 ;
  wire  \inst_doa_mux_b29/B0_2 ;
  wire  \inst_doa_mux_b29/B0_3 ;
  wire  \inst_doa_mux_b29/B1_0 ;
  wire  \inst_doa_mux_b29/B1_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b3/B0_2 ;
  wire  \inst_doa_mux_b3/B0_3 ;
  wire  \inst_doa_mux_b3/B1_0 ;
  wire  \inst_doa_mux_b3/B1_1 ;
  wire  \inst_doa_mux_b30/B0_0 ;
  wire  \inst_doa_mux_b30/B0_1 ;
  wire  \inst_doa_mux_b30/B0_2 ;
  wire  \inst_doa_mux_b30/B0_3 ;
  wire  \inst_doa_mux_b30/B1_0 ;
  wire  \inst_doa_mux_b30/B1_1 ;
  wire  \inst_doa_mux_b31/B0_0 ;
  wire  \inst_doa_mux_b31/B0_1 ;
  wire  \inst_doa_mux_b31/B0_2 ;
  wire  \inst_doa_mux_b31/B0_3 ;
  wire  \inst_doa_mux_b31/B1_0 ;
  wire  \inst_doa_mux_b31/B1_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b4/B0_2 ;
  wire  \inst_doa_mux_b4/B0_3 ;
  wire  \inst_doa_mux_b4/B1_0 ;
  wire  \inst_doa_mux_b4/B1_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b5/B0_2 ;
  wire  \inst_doa_mux_b5/B0_3 ;
  wire  \inst_doa_mux_b5/B1_0 ;
  wire  \inst_doa_mux_b5/B1_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b6/B0_2 ;
  wire  \inst_doa_mux_b6/B0_3 ;
  wire  \inst_doa_mux_b6/B1_0 ;
  wire  \inst_doa_mux_b6/B1_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b7/B0_2 ;
  wire  \inst_doa_mux_b7/B0_3 ;
  wire  \inst_doa_mux_b7/B1_0 ;
  wire  \inst_doa_mux_b7/B1_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b8/B0_2 ;
  wire  \inst_doa_mux_b8/B0_3 ;
  wire  \inst_doa_mux_b8/B1_0 ;
  wire  \inst_doa_mux_b8/B1_1 ;
  wire  \inst_doa_mux_b9/B0_0 ;
  wire  \inst_doa_mux_b9/B0_1 ;
  wire  \inst_doa_mux_b9/B0_2 ;
  wire  \inst_doa_mux_b9/B0_3 ;
  wire  \inst_doa_mux_b9/B1_0 ;
  wire  \inst_doa_mux_b9/B1_1 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i0_012;
  wire inst_doa_i0_013;
  wire inst_doa_i0_014;
  wire inst_doa_i0_015;
  wire inst_doa_i0_016;
  wire inst_doa_i0_017;
  wire inst_doa_i0_018;
  wire inst_doa_i0_019;
  wire inst_doa_i0_020;
  wire inst_doa_i0_021;
  wire inst_doa_i0_022;
  wire inst_doa_i0_023;
  wire inst_doa_i0_024;
  wire inst_doa_i0_025;
  wire inst_doa_i0_026;
  wire inst_doa_i0_027;
  wire inst_doa_i0_028;
  wire inst_doa_i0_029;
  wire inst_doa_i0_030;
  wire inst_doa_i0_031;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i1_009;
  wire inst_doa_i1_010;
  wire inst_doa_i1_011;
  wire inst_doa_i1_012;
  wire inst_doa_i1_013;
  wire inst_doa_i1_014;
  wire inst_doa_i1_015;
  wire inst_doa_i1_016;
  wire inst_doa_i1_017;
  wire inst_doa_i1_018;
  wire inst_doa_i1_019;
  wire inst_doa_i1_020;
  wire inst_doa_i1_021;
  wire inst_doa_i1_022;
  wire inst_doa_i1_023;
  wire inst_doa_i1_024;
  wire inst_doa_i1_025;
  wire inst_doa_i1_026;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i2_009;
  wire inst_doa_i2_010;
  wire inst_doa_i2_011;
  wire inst_doa_i2_012;
  wire inst_doa_i2_013;
  wire inst_doa_i2_014;
  wire inst_doa_i2_015;
  wire inst_doa_i2_016;
  wire inst_doa_i2_017;
  wire inst_doa_i2_018;
  wire inst_doa_i2_019;
  wire inst_doa_i2_020;
  wire inst_doa_i2_021;
  wire inst_doa_i2_022;
  wire inst_doa_i2_023;
  wire inst_doa_i2_024;
  wire inst_doa_i2_025;
  wire inst_doa_i2_026;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;
  wire inst_doa_i3_009;
  wire inst_doa_i3_010;
  wire inst_doa_i3_011;
  wire inst_doa_i3_012;
  wire inst_doa_i3_013;
  wire inst_doa_i3_014;
  wire inst_doa_i3_015;
  wire inst_doa_i3_016;
  wire inst_doa_i3_017;
  wire inst_doa_i3_018;
  wire inst_doa_i3_019;
  wire inst_doa_i3_020;
  wire inst_doa_i3_021;
  wire inst_doa_i3_022;
  wire inst_doa_i3_023;
  wire inst_doa_i3_024;
  wire inst_doa_i3_025;
  wire inst_doa_i3_026;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i4_003;
  wire inst_doa_i4_004;
  wire inst_doa_i4_005;
  wire inst_doa_i4_006;
  wire inst_doa_i4_007;
  wire inst_doa_i4_008;
  wire inst_doa_i4_009;
  wire inst_doa_i4_010;
  wire inst_doa_i4_011;
  wire inst_doa_i4_012;
  wire inst_doa_i4_013;
  wire inst_doa_i4_014;
  wire inst_doa_i4_015;
  wire inst_doa_i4_016;
  wire inst_doa_i4_017;
  wire inst_doa_i4_018;
  wire inst_doa_i4_019;
  wire inst_doa_i4_020;
  wire inst_doa_i4_021;
  wire inst_doa_i4_022;
  wire inst_doa_i4_023;
  wire inst_doa_i4_024;
  wire inst_doa_i4_025;
  wire inst_doa_i4_026;
  wire inst_doa_i5_000;
  wire inst_doa_i5_001;
  wire inst_doa_i5_002;
  wire inst_doa_i5_003;
  wire inst_doa_i5_004;
  wire inst_doa_i5_005;
  wire inst_doa_i5_006;
  wire inst_doa_i5_007;
  wire inst_doa_i5_008;
  wire inst_doa_i5_009;
  wire inst_doa_i5_010;
  wire inst_doa_i5_011;
  wire inst_doa_i5_012;
  wire inst_doa_i5_013;
  wire inst_doa_i5_014;
  wire inst_doa_i5_015;
  wire inst_doa_i5_016;
  wire inst_doa_i5_017;
  wire inst_doa_i5_018;
  wire inst_doa_i5_019;
  wire inst_doa_i5_020;
  wire inst_doa_i5_021;
  wire inst_doa_i5_022;
  wire inst_doa_i5_023;
  wire inst_doa_i5_024;
  wire inst_doa_i5_025;
  wire inst_doa_i5_026;
  wire inst_doa_i6_000;
  wire inst_doa_i6_001;
  wire inst_doa_i6_002;
  wire inst_doa_i6_003;
  wire inst_doa_i6_004;
  wire inst_doa_i6_005;
  wire inst_doa_i6_006;
  wire inst_doa_i6_007;
  wire inst_doa_i6_008;
  wire inst_doa_i7_000;
  wire inst_doa_i7_001;
  wire inst_doa_i7_002;
  wire inst_doa_i7_003;
  wire inst_doa_i7_004;
  wire inst_doa_i7_005;
  wire inst_doa_i7_006;
  wire inst_doa_i7_007;
  wire inst_doa_i7_008;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[10]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  reg_sr_as_w1 addra_pipe_b2 (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[2]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00000000000000000000000000000000000000000000000152935E03E6666666),
    .INITP_01(256'h000000000000000000000000000000000000000000B333333430049600000003),
    .INITP_02(256'hFB02C75F4BEB2BE8205EE9A1C94094599321CA38000000000000000000000000),
    .INITP_03(256'hA18614AACAB40DE1CCCCCCC5681AE20287D3985250AC972C79B43213AE97F3D7),
    .INIT_00(256'h3793139313931393139313931393139313931393139313931393139313931393),
    .INIT_01(256'h670B670B73EF13E31313238313179313E3132393971393736F0B232323231313),
    .INIT_02(256'h000000000000000000000000000000000000000000000000000000000000670B),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h2323232323232323232323232323232323232323232323232323238B238B0B13),
    .INIT_09(256'h83038303830B830B830B03038313172383131723630313170BEFEF8BEF138B23),
    .INIT_0A(256'h000000000000000B138B83038303830383038303830383038303830383038303),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h9402788484010000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h000000000000000000000000000000000000000000002CB4B40A30A4A4052094),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h931393B7B7EF13931393B7B7EFEF2313B737EF23136F1383EF231303B7670000),
    .INIT_14(256'h13376723B76FEF13EF1313B723233723136FEF13EF13372323136F131383EF13),
    .INIT_15(256'h23231367232323136703E3131393936733B30363336393939313036F23676383),
    .INIT_16(256'h6713038313239393B3B3139313B71313639313838323B3831383836383EF2313),
    .INIT_17(256'h131333831393B70363EF23132323136F131383EF231393136F136FB393139313),
    .INIT_18(256'h939393B793B3936713038313233393B73313939363139393B393030323838333),
    .INIT_19(256'h23131337936FEF13936713038303038363EF13931393A323232323136F23B333),
    .INIT_1A(256'h03333393EF1323231363936F131383E393232313933793B7EF231367131383EF),
    .INIT_1B(256'h136723236303B39313B76393676F1333938303B393EF132323136393676F1383),
    .INIT_1C(256'h03830383130383E31393E7138363836393B39393131313232323232337231367),
    .INIT_1D(256'h8303830383038303830383038303830383038303830383038303838303036713),
    .INIT_1E(256'h03B7672313233723376303B76F9323672323232393B763139313371313136713),
    .INIT_1F(256'h3767130383736383B76313236303B7EF132323136F136723B723132337233763),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_008,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000058080000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000002210000000000),
    .INITP_02(256'hEC4010BF03FFE694016E7F9A1410420038760090000000000000000000000000),
    .INITP_03(256'h831D0955956EFB4E000000000025C000372190202041FE001400400BFE07FFC3),
    .INIT_00(256'h2007070707060606060505050504040404030303030202020201010101000000),
    .INIT_01(256'h40B240B2001002A48203901303030202FE8290C20A0200000030939291908080),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000004062),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h969594939291909796959493929190979695949392919097969591A090205080),
    .INIT_09(256'h92929191915090509090925012020A5012020A108414020AE010006210009097),
    .INIT_0A(256'h000000000000000080A097979797969696969595959594949494939393939292),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0100000101000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000010100000101000001),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'hC203430A2B0002C203430A2B00F8D6820BC2089380088090F89380D20B400000),
    .INIT_14(256'h820340D203F818021842022A93910A9280F8180218022A939280008002900002),
    .INIT_15(256'h979680408A90913B400A8302BBFBAB4082C30AF442C7ABEB8B8393F89240CAA3),
    .INIT_16(256'h408092900211EBCBF3FB8B43A383BBEB8943EB0B13C0C313EB9213C20BF89382),
    .INIT_17(256'hAB8BBB13ABC3431386F8938297968008800290F893020280F802F8F3EB8BCB83),
    .INIT_18(256'hCB43EB83CBFBC3408092900211BBC383B3BBE3BBCE03EBCBFBAB0B13C092A3C3),
    .INIT_19(256'h9382802A82F808020240809492A2929088F802820202839794959680F811B3BB),
    .INIT_1A(256'h9232CA030082939280E50300800290CDC3D1D083C30BC30B0093804080029010),
    .INIT_1B(256'h0240D1D0C5D2C3C38A0BE203400080FAE39092CB030082939280E60340008090),
    .INIT_1C(256'h959494928292904E0242C04212C413C6FB2B040202C58497929394950A968040),
    .INIT_1D(256'h9797979796969696959595959494949493939393929292929191919091904080),
    .INIT_1E(256'hD30B40D003910B920B8BD30BF8C3D04012101211C34308838302E3843B030080),
    .INIT_1F(256'h2A4080929000C2D30B0D3AD780D30BF882939280F80240D70BD003910B920B8B),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_017,inst_doa_i0_016,inst_doa_i0_015,inst_doa_i0_014,inst_doa_i0_013,inst_doa_i0_012,inst_doa_i0_011,inst_doa_i0_010,inst_doa_i0_009}));
  // address_offset=0;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000001500984200000000),
    .INITP_01(256'h0000000000000000000000000000000000000000013FFFC000022169FFFE0000),
    .INITP_02(256'h048217A00014C000212000110600D86224482CA0000000000000000000000000),
    .INITP_03(256'h01001C5495280128FFFF00000100080201048040009512216680201810014400),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h00810081040000AD11113D0181007000A9110121FF700004208000000000C000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'hF8F4F0ECE8E4E05C5854504C484440BCB8B4B0ACA8A4A01C1814040004008000),
    .INIT_09(256'h9080706050801080008100010101FF090151FF01820181FF00A4C400340080FC),
    .INIT_0A(256'h00000000000000000000F0E0D0C0B0A090807060504030201000F0E0D0C0B0A0),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h2100D10000A0003100A1000020C3A98100000404C0A440307304C0E100000000),
    .INIT_14(256'h0580002980C764016071E10004240020C0C724402001000420C0F04004303004),
    .INIT_15(256'h04208000312D01F10021BD00050541003D3521353D354545410111B73D0001FD),
    .INIT_16(256'h00806070043D3D3D393541FD05FF054135FD4521112D39014530112921372C01),
    .INIT_17(256'h4141350105FD001181F72C01042080C440C030170400FCC0570057393D453D05),
    .INIT_18(256'h050541FF4135050080607004393D05FF3DF90505B1FD4141350521113D300139),
    .INIT_19(256'h04E1C00001272401FC008040503C6070A537003CC004000448242080173D3D35),
    .INIT_1A(256'h20292104F0010420C0A97C8040FC30B5210139B1010001003004C000400030D4),
    .INIT_1B(256'h0000312D010129010D00A97C00A04029FD3020210400010420C0A97C00A04030),
    .INIT_1C(256'h203040500260704D21050101110101010526800001010104504C482400208000),
    .INIT_1D(256'hF0E0D0C0B0A090807060504030201000F0E0D0C0B0A090807060501000010080),
    .INIT_1E(256'h01000039042D002900010100671139003D41AD350100BDBD0101AB01F1110000),
    .INIT_1F(256'h00004020300001010001098181F100C3010420C013FC00B90039042D00290001),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_026,inst_doa_i0_025,inst_doa_i0_024,inst_doa_i0_023,inst_doa_i0_022,inst_doa_i0_021,inst_doa_i0_020,inst_doa_i0_019,inst_doa_i0_018}));
  // address_offset=0;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000004508980200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000008000000006630400000001),
    .INIT_02(256'h044307A000144014212000110460F44285012C20000000000000000000000000),
    .INIT_03(256'h000014000008F969000000000100000200048040008510A06680201810014400),
    .INIT_04(256'h00BD00221000040004020001E041294000089000292500002060367000040C11),
    .INIT_05(256'h000080198000000894492060807FFE000220003FFE5319A500033081A000000D),
    .INIT_06(256'h80400000D2120448080000131A41C0600040B650008000D405C8022100004000),
    .INIT_07(256'h36AF40400000006619002040206008010620200098400800240010000185C861),
    .INIT_08(256'h00D0104002000008100642A40002008204061800010000400551010818200440),
    .INIT_09(256'h02000003100041009000C880000020400002140F0C00008B0060C0182008060A),
    .INIT_0A(256'h08A04880008000008201000000050182048000401284002E00A40828400201A0),
    .INIT_0B(256'h00808342000016EDB3500140491531000001080040A00018140024A544000000),
    .INIT_0C(256'h0041080017F0902D840080280A02D800D80400021000E12440082202080000C0),
    .INIT_0D(256'h46184D00324A0000001001060000802802200C080400800160D0446840090405),
    .INIT_0E(256'hC920E04020200A0007060220000600010088001C008941009215480000610682),
    .INIT_0F(256'h46000880E00A4302621900424004408002040006000108100240280100800A40),
    .INIT_10(256'h8843000200018041044020000001900000001101901000824204001080204080),
    .INIT_11(256'h410810010004400804008090100440028004068000500800840180204000A054),
    .INIT_12(256'h03180400740620020090481020008DC85500020401A90400812108A000000821),
    .INIT_13(256'h870150346C743641D430CE0C0A8482500745042810804B184D00500400000407),
    .INIT_14(256'h0000000000001400112522509117CC820092015AFF02008A2175F60A8082ED06),
    .INIT_15(256'h0A843235A7001000649249249249249240887002070000000408420009000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_027 (
    .addra(addra),
    .clka(clka),
    .dia({open_n195,open_n196,open_n197,open_n198,open_n199,open_n200,open_n201,1'b0,open_n202}),
    .rsta(rsta),
    .doa({open_n217,open_n218,open_n219,open_n220,open_n221,open_n222,open_n223,open_n224,inst_doa_i0_027}));
  // address_offset=0;data_offset=28;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000100880200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000002212000000001),
    .INIT_02(256'h040311A0001440042120001104A0D862850E0CB0000000000000000000000000),
    .INIT_03(256'h01151D549528F06800000000010008020104804000850A202680401810014400),
    .INIT_04(256'h80B900223000040008020001A0412940000A9000212500088060B23000042C1B),
    .INIT_05(256'h4000001B810000089441006AA10002020320504000C1108C000010003000000D),
    .INIT_06(256'h80C00000D0022411A0000400001401000040B440009100540560026B40004204),
    .INIT_07(256'h260940C8804001768000006000C284200E6640009A400800040004000901C841),
    .INIT_08(256'h00D21660828A5089110D4240012E0180040C38800B250180050002887AE7255E),
    .INIT_09(256'h02000003300041002000EEC009002040000214340C4D908B0060C01820080602),
    .INIT_0A(256'h0DA8488000A810008001000000050092048010C01A84002C00200800400001A0),
    .INIT_0B(256'h00000042100014A9225010084D10910002010D0840A00014840026A424000401),
    .INIT_0C(256'h1041080017F0006D840080000A10D048D09400021000E12440082212080080C0),
    .INIT_0D(256'h46084D00324A0000001001060000802802200C080400800160D0446840090405),
    .INIT_0E(256'h0920000028200E0807060220000600010080001C02894900D011480000000682),
    .INIT_0F(256'h46000880E0024388621D0043400040000204000600010C500240000000081108),
    .INIT_10(256'h8843040200018000001020080000100002001901901000000280069AD2B04080),
    .INIT_11(256'h4908110100044008040080901004C0028004040480500200042580250220A044),
    .INIT_12(256'h071804007406000A209048102050EDCC15000B0401A90400810008A004028CA3),
    .INIT_13(256'h048606428A02C11600C6819302D001400644000010804B184D06508000000404),
    .INIT_14(256'h000000000018C0211004208420000227500040000052570080780011041000A0),
    .INIT_15(256'h307209C000020000000000000000000000618000AD000000019A8296A0000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_028 (
    .addra(addra),
    .clka(clka),
    .dia({open_n256,open_n257,open_n258,open_n259,open_n260,open_n261,open_n262,1'b0,open_n263}),
    .rsta(rsta),
    .doa({open_n278,open_n279,open_n280,open_n281,open_n282,open_n283,open_n284,open_n285,inst_doa_i0_028}));
  // address_offset=0;data_offset=29;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000100880200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000002214C00000001),
    .INIT_02(256'h044215A000144004212000110660F462244D28A0000000000000000000000000),
    .INIT_03(256'h000014000008F148000000000100000200008444089500A16680601810014400),
    .INIT_04(256'h80B900223000042008020801A041284000028000216500002060B67000042C1B),
    .INIT_05(256'hC0A0001B0100000000000062800002020000004000E191AD000230011000000D),
    .INIT_06(256'h80C00000D2122441A00000010A0000000040B250018040D705EC026B40004006),
    .INIT_07(256'h260940C800400174A903006020A28CB3462000009AC00800240000000105C861),
    .INIT_08(256'h10C2144002000089110D4240012A0100008828808F7581C0054103983AE7255E),
    .INIT_09(256'h0200000310004110B60CEC001904200000021404AC48108B0000C00020080E0A),
    .INIT_0A(256'h0DA04880008010008201000010050000048004C21A54080E00A40808400001A0),
    .INIT_0B(256'h10800042100014A92250000049143100020004A808B00018100036A564000401),
    .INIT_0C(256'h1041080017F0006D840080000A00D000D00400021000E12440082212080080C0),
    .INIT_0D(256'h46084D00324A0000001001060000803802200C080400800160D0446840090405),
    .INIT_0E(256'h0920A00028200E0807970220000600010080001C00014900C011482209000682),
    .INIT_0F(256'h46000880E002430062190042401448A00200008680030C500240280000081108),
    .INIT_10(256'h88430402000180010400200000001000020010019000802242048412C0B04080),
    .INIT_11(256'h4908010100040008040008804004C0000200040080502A008425802D0220A044),
    .INIT_12(256'h071804007406000A20904810200089C81400022001A90400812908A004000823),
    .INIT_13(256'h858D76F6EEF6F33FD5F6CFBF6F56C1590D45242810804B184D06508000000404),
    .INIT_14(256'h000000000078D4A155F7F2F9B773DFB7FDB6DB3FFF7FFFA79B7DFEFFAFBEFCFE),
    .INIT_15(256'h27FFFFF7FF000002000000000000000004FFF002AD00000007FEFEDF44000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_029 (
    .addra(addra),
    .clka(clka),
    .dia({open_n317,open_n318,open_n319,open_n320,open_n321,open_n322,open_n323,1'b0,open_n324}),
    .rsta(rsta),
    .doa({open_n339,open_n340,open_n341,open_n342,open_n343,open_n344,open_n345,open_n346,inst_doa_i0_029}));
  // address_offset=0;data_offset=30;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000000000000000050A8C0200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000006630000000001),
    .INIT_02(256'h044351A0001440042120C8110440D440204508A0000000000000000000000000),
    .INIT_03(256'h000014000008F168000000000100000200008040008510216480481810014400),
    .INIT_04(256'h80BD0026B400042008020001A0412940000A9000212100000060323000040C13),
    .INIT_05(256'h0000801A4000401000080862800002000260004000E1908C000230813000000D),
    .INIT_06(256'h80C00000D0022401A00000000000001000403000008000540560026B40004000),
    .INIT_07(256'h2609404080C000663000204020000400062220009AC40800040000000185C861),
    .INIT_08(256'h1052144822000008100442240002002004020800811000080541081018202542),
    .INIT_09(256'h02000103300041101404EC00090024800A02140DCC25008B0060C01820080808),
    .INIT_0A(256'h0408408000C0500080A1000000050192048014421AD4080E00A40828400201A0),
    .INIT_0B(256'h000004420000102100500000491431000215040040A00010040034A504000415),
    .INIT_0C(256'h10410C121FF0006D8420A0000A02D008D01400031000F1346008A312088080C0),
    .INIT_0D(256'hC6084D00324A0000015003060000803812200C882440940160D0C46860090405),
    .INIT_0E(256'hCD60800028200A0005D32220480600000089009C02814900C011482000000682),
    .INIT_0F(256'h46880080E00561C0660DAF404004408002000006000108100240000080480148),
    .INIT_10(256'h80420200000DCAC000502810000110000000190192B0A0A24A048C52C0B16000),
    .INIT_11(256'h4908110100044008040028844014C0000000040180500000042580204240A010),
    .INIT_12(256'h071804007406001F21BA489020008DC85D00022001A90400812908B004000821),
    .INIT_13(256'h838776F6EEF6F337D5F6DA956F4403100741040411804F184D06D08000002404),
    .INIT_14(256'h0000000000631421152162DDB0001E300192C800005F57229B60009B282000F4),
    .INIT_15(256'h1FFBFFF6F8020000000000000000000004F78002A200000005F0D217A1000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_030 (
    .addra(addra),
    .clka(clka),
    .dia({open_n378,open_n379,open_n380,open_n381,open_n382,open_n383,open_n384,1'b0,open_n385}),
    .rsta(rsta),
    .doa({open_n400,open_n401,open_n402,open_n403,open_n404,open_n405,open_n406,open_n407,inst_doa_i0_030}));
  // address_offset=0;data_offset=31;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000100880200000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000006630000000001),
    .INIT_02(256'h044211A000144004212000110460C440A14408A0000000000000000000000000),
    .INIT_03(256'h00011C000008F968000000000100080201008040008512206480401810014400),
    .INIT_04(256'h00AC0026B400042008020001A0412940000A9000212100000060323000040C13),
    .INIT_05(256'h8000001A000000000000206AA00002020040000000C111AD000010802000000D),
    .INIT_06(256'h80C0000050022401A0000000000000000040B000008000540560026B40004200),
    .INIT_07(256'h26094040804000641101204000000410440000009A400000000000000185C861),
    .INIT_08(256'h0040104822000008100442240002000004030810811000000541001858202542),
    .INIT_09(256'h02000003910041000404EE4000002040000214046801008B0000C00020080000),
    .INIT_0A(256'h0C80488000C0400080A1000000050092048004421A40080E00A40808400001A0),
    .INIT_0B(256'h0000004200001225815011484D14910002010C8048B00018100036A524000401),
    .INIT_0C(256'h1041080017F0006D840080000A02D008D01400021000E12440082212080080C0),
    .INIT_0D(256'h46084D00324A0000001001060000803802200C080400800160D0446840090405),
    .INIT_0E(256'h0920A00028200E0807972220400600010088001C02814900C011482000000682),
    .INIT_0F(256'h46000088F0804182620D00404004408002040086800308100240000000080108),
    .INIT_10(256'h884306000005C0410410200000011080020019019010A08242048412C0B04000),
    .INIT_11(256'h4908152100044008040088905004C00282040404805028008425802C0220A044),
    .INIT_12(256'h071804007406000A2090481020008DCC5500026401A90400812908A004000A23),
    .INIT_13(256'h000000000000000000000000035601580755240210804B184D06508000000404),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_031 (
    .addra(addra),
    .clka(clka),
    .dia({open_n439,open_n440,open_n441,open_n442,open_n443,open_n444,open_n445,1'b0,open_n446}),
    .rsta(rsta),
    .doa({open_n461,open_n462,open_n463,open_n464,open_n465,open_n466,open_n467,open_n468,inst_doa_i0_031}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h600AC0C139BCC1DEB04D5003280142AEA71389A032331B0B407622B70C058E83),
    .INITP_01(256'h04D50034CE1C79EAD6F55283CDE660C5E5836A8001974E0E6E61C572C1B54018),
    .INITP_02(256'h780B4CC36719956E4224EB28C62E368D00562331B0D680E98A5624939BCC1DEB),
    .INITP_03(256'h54132A992E040959DC51916E13A7189917BBBB986074F46262F60760036A310C),
    .INIT_00(256'h83038363B737932323232303231367131383EF2313133767138363EFEF231313),
    .INIT_01(256'h03B7EF23232323232313133767131383EF23136F03EF136383EF139367138303),
    .INIT_02(256'h232313836323836F13EF139363EF13931383671313038303830383638337B737),
    .INIT_03(256'h130393036713830383038313EF639303836393EF131363138363139313232323),
    .INIT_04(256'h6FEF1367138303836313B7132323231367136F136F2313EF13E3932333031363),
    .INIT_05(256'h93EF1337EFEF2323239313231393133737932313EF2323232323232323231313),
    .INIT_06(256'hEF63938303EF83B393671313830383038303830383E363831393EF9313B737B7),
    .INIT_07(256'hEF139313630313136F136FEF13EF13EF13931363031313638303931303EF6F13),
    .INIT_08(256'h1337EFEF2323239393231393133737932313EF232323232323232313136F136F),
    .INIT_09(256'h03B3936713130383038303830383EF133793EFE363839313EF931337B73713EF),
    .INIT_0A(256'h2323232323232313136FEF1363931383EF931393130383EF6F93EF63938303EF),
    .INIT_0B(256'h13B737B73713EF1337EFEF2323239393231393133737932313EF232323232323),
    .INIT_0C(256'h8303EF03B39367131383038303830383038303830383E3638337B7379313EF93),
    .INIT_0D(256'h131363136313136393131383EF9313138303EF13EF23131393936F93EF639393),
    .INIT_0E(256'h13B39303038383EF23232313933393B39333B30383036303139383EF13631363),
    .INIT_0F(256'hEFEF2323239313231393133737932313EF23232323232323232313136F136FEF),
    .INIT_10(256'h03EF83B393671313830383038303830383E363831393EF9313B737B793EF1337),
    .INIT_11(256'h93136303936F936FEF13EF13EF139313630393631303931383EF6F13EF639383),
    .INIT_12(256'h13038303830383EF1337638337B73703B7EF2323232323231313376F936FEF13),
    .INIT_13(256'h13232323232323232313671367131383EF23136F13EF139363EF139313836713),
    .INIT_14(256'h13931363EF13931303633783B783B763636383B393131363136363B3831393B3),
    .INIT_15(256'h6F136F136F63936363638313131393131313939313EF139313638363833363EF),
    .INIT_16(256'hEF1337E3EF131383B713EF1337636F9313236F936F13EF9323133763130393E3),
    .INIT_17(256'h6F139313936363836FE363638323139363136367130383038303830383E79313),
    .INIT_18(256'h232323230323B7136F139363836F936FE36F1393E3636383236FE393931323E3),
    .INIT_19(256'hEF139313036F13831303839313830383038303636383B737B793139323232323),
    .INIT_1A(256'h6F1393E3E3836F13EF13939363B3630313931393EF136363EF13931313EF1363),
    .INIT_1B(256'h2313233723139337B7239337B7239337B7239337B76713830383038303830383),
    .INIT_1C(256'h0383EF136323938303EF931393B70313EF2323139313931393932313B7371393),
    .INIT_1D(256'h93B7EF1393B763EF6713831303832393B7639393233723832313836713130383),
    .INIT_1E(256'hEF37B737B73737B7EFEF232323932323232323238323230323136F93B76FEF13),
    .INIT_1F(256'h6313E3132313E3136F936313E3931313236F136313630393836F231383639393),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_008,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=1024;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h44AC8806E700002718038000802029FA800E104009200006801011000C000210),
    .INITP_01(256'h8038000A800F020DA98120AE3000007278C01C00005E09B98000809C600E0005),
    .INITP_02(256'hFDAF2000208BE0BCA120001C8634E06000009200004D003D1764406E70000271),
    .INITP_03(256'h3A0AC660FF64082C450351000704041C4AEEE800FF5F000028000F000897F9FF),
    .INIT_00(256'h929290082C2C829793949592968040800290109382802A40809088F810938280),
    .INIT_01(256'hD20B1095979293949682802A40800290109380F81210C2C31310820240809494),
    .INIT_02(256'h959680E3C3D4D3F802100242841842C2031240800295949492929032932D2C0C),
    .INIT_03(256'hC41203534080949492929002F8C2FB63238E83F804C20B04D4C702C282939497),
    .INIT_04(256'hF8104240809292900E022A02939192804002F802F85402F842C8C3900354CBC4),
    .INIT_05(256'h0410822AF8109794960385858202032A2B039382109091929394959697930280),
    .INIT_06(256'hF8C4FB63A3F8D2038B408002959595959494929290C9A6930484F882C22D2D2D),
    .INIT_07(256'h104202030E130403F804F810C2F802108202030A130403006B6B434253F8F884),
    .INIT_08(256'h822AF8109794960384858202032A2B0393821095969091929394970280F804F8),
    .INIT_09(256'hD2C34B408002959595949492929010822A82008962930284F882822D2D2D0410),
    .INIT_0A(256'h979091929394970280F81042CAFB822310020303021313F8F842F8C4FB23A3F8),
    .INIT_0B(256'h822D2D2D2D0410822AF8109196900384878202032A2B03958210939495969596),
    .INIT_0C(256'h23A3F8D2C34B408002969696969595959594949292908E62932E2E2E0284F882),
    .INIT_0D(256'hC203C702C14203C4FB820323100203029323F8C2189182034203F842F8C4FB86),
    .INIT_0E(256'h42C28393939312189192938A02424B438BC2C613131381A3C203161082CB03C4),
    .INIT_0F(256'hF8109794960385858202032A2B039382109091929394959697930280F882F810),
    .INIT_10(256'hA3F8D2038B408002959595959494929290C9A6930484F882C22D2D2D0410822A),
    .INIT_11(256'h02030E1303F8C3F810C2F802108202030A130307036B434253F8F884F8C4FB63),
    .INIT_12(256'h0295949492929010822A35932D2C0CD20B1095979293949682802AF8C3F81042),
    .INIT_13(256'h82909192939495979680400240800290F89380F8021002428C1842C203124080),
    .INIT_14(256'h0202838818028203D5FB2DD50BD40B8EC1C2E3030303044302C6C7C223030382),
    .INIT_15(256'hF884F8020081038ECBC2E20703010404030203838418820203C3D4C823058B18),
    .INIT_16(256'h08822A8C108442922A8210822A8BF8C383C0F8C400021002C0822A8DBBE30389),
    .INIT_17(256'hF883C383C34BCCE7F88BB3C4E25083C3C882B940809595959494929290C08202),
    .INIT_18(256'h95979091D5960B80F80202CCA3F8C3F8B5F883C383C5C6E250F8B043C383C0BE),
    .INIT_19(256'h180282031208809242949482C39595959590928430532D2D0D04048292939394),
    .INIT_1A(256'hF883C30E47A3F80508C202C4EAC309E3038304841002CD881842028302184288),
    .INIT_1B(256'h9182920B9380C30B2B94C30B2B95C30B2B96C30B2B4080959595959494929290),
    .INIT_1C(256'h929010028B81F3A31300C203032A128410909302C2030304030412832A130203),
    .INIT_1D(256'hC22A1002C22A82F8408092429290C6C30BCA02FB930A91E39280134080029492),
    .INIT_1E(256'hF02E2D2D2C2C2D2D08F8819191F3929394959697A39093139280F8C22AF81042),
    .INIT_1F(256'h8A037ABBD0838F0300064C037403BB43D0F8038B038ED30313F8D003138D8203),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_017,inst_doa_i1_016,inst_doa_i1_015,inst_doa_i1_014,inst_doa_i1_013,inst_doa_i1_012,inst_doa_i1_011,inst_doa_i1_010,inst_doa_i1_009}));
  // address_offset=1024;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hC0888120342FFC20480207FCE0412040000A9000282500088060367000042C09),
    .INITP_01(256'hC000FFC18000021890002B42807FFF020140003FFE53180C0BFD188120283FE4),
    .INITP_02(256'h80008800D0040E490D9004401814C16000402400009100530464020302FFC204),
    .INITP_03(256'h522748C8000001660903006020E288314E6660009A40090104001C000904C061),
    .INIT_00(256'h506070A5000001044C482401208000400030040401C0000040300167A40481C0),
    .INIT_01(256'h6100042404504C4820718000004000305404C00701346225017452B100803040),
    .INIT_02(256'h24208021010131B72174D20101B401C20801008000203040506070BD52000000),
    .INIT_03(256'h01010011008030405060700097B9FD21F18201E70402010001810001014C4804),
    .INIT_04(256'h77F4E1004010203001FD0024042420C00000A700A749014701C90521393109A2),
    .INIT_05(256'h00F4A100573400503C20803C1120F1000014281104C8A4A05C5854504C841440),
    .INIT_06(256'hD739FDF15007013E0A00C00030405060708090A0B082BE700001473002000000),
    .INIT_07(256'hE0722020310100014706B790420701D0122020B1010001315159D12121A77706),
    .INIT_08(256'h91003710004C3C20803CF120D10000282811E424205854504C48042880870607),
    .INIT_09(256'h013E090080000010203040506070C0F1000194823D70000127300200000000D0),
    .INIT_0A(256'h5CD8D4D0CCC88404000780B2010582F5E02020D12261714737057739FDF150A7),
    .INIT_0B(256'h020000000000408100A780804CBC20A03C7120510000042811506C686460A4A0),
    .INIT_0C(256'hF170D7013E0900000030405060708090A0B0C0D0E0F0023D9000000000018750),
    .INIT_0D(256'h42100113B9E308B93DB304A1A020208210A5F703B03420E001D127059739FD01),
    .INIT_0E(256'hA22F01102030413030383C0901290D29052B33D19181BD01038C719072390C39),
    .INIT_0F(256'h17F000503C20803C7120410000082811C0C8A4A05C5854504C840840570537D0),
    .INIT_10(256'h50C3013E0A00C00030405060708090A0B082BE70000107300200000000B0E100),
    .INIT_11(256'h20203101004705C76042D301A0422020B10100BD0141D121216377069339FDF1),
    .INIT_12(256'h00203040506070504100BD520000006100F02404504C4820218000870527C082),
    .INIT_13(256'h01D8D4D0CCC8A484A0000004004000308704C0872130B2190170019218010080),
    .INIT_14(256'h1A0102012002921802D60051006100A63539014924800081003935210124802D),
    .INIT_15(256'hD7066705B0BD2025C5410170882024800000010000200000808212811A4A81D0),
    .INIT_16(256'hE44100A22012B102008080C1009947050501972280FC4001014100817D010102),
    .INIT_17(256'h4705050505337105A78125B1013D0505B105A500008090A0B0C0D0E0F0020020),
    .INIT_18(256'h544CC8A461500040E70000010107056725A70505A54541013D07251105050125),
    .INIT_19(256'hE00192180270C090018070020230405060B0A0023E52000000000001A0845C58),
    .INIT_1A(256'h170505350101172264D201014D49810101020101B40102016001010119400181),
    .INIT_1B(256'h240120003DC0F100003DF100003D8100003DC1000000C030405060708090A0B0),
    .INIT_1C(256'h2030900102BD09912024C10000002001D0480401A161001800283C0100000130),
    .INIT_1D(256'h210024E1E10081C700401001203081010081E1090400249120C0200040000010),
    .INIT_1E(256'h570000000000000064F7BD64A405605C5854504C91C88420A040770100072401),
    .INIT_1F(256'hB91039FD81FD31082000B924B9F4FDFD817708396CB581042097B904203D016C),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_026,inst_doa_i1_025,inst_doa_i1_024,inst_doa_i1_023,inst_doa_i1_022,inst_doa_i1_021,inst_doa_i1_020,inst_doa_i1_019,inst_doa_i1_018}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00C8997442C52B9F3F79B4495B6BB75D5160EBA53A2D77B6632A74C4945DDA75),
    .INITP_01(256'h241B1412567081692661892624A838930A02C5800A499AA228008A002AAA27F6),
    .INITP_02(256'h5256964B9895A000B1496044A045702C051B0258152B1514B1280B1258081141),
    .INITP_03(256'hCC034090D40315695A5606A0526253D9859E5256962973132800210894E5699E),
    .INIT_00(256'h93EFEF13E3838393EF136F938303EF138333E30303E3136F23938303EF13E383),
    .INIT_01(256'h232313131313131303E303631363136F23231313EF1383EF139313EFEF136393),
    .INIT_02(256'h6FA3B30383EF136F93EF13E383838383EFB39383A333031383EF33B333139363),
    .INIT_03(256'h03236313836F2323EF13931383EFEFEF138303EF13639383836393EF63136313),
    .INIT_04(256'h23139313138303836383838383EF13B393631303A3338383EF3333B313936303),
    .INIT_05(256'h672333130393130367131303836FEF1393E39383A3336F93EF136F2323E39323),
    .INIT_06(256'h23B7EF132323136703B7676723B723B76723B723B7671303836723B393831303),
    .INIT_07(256'h133313EF932323239313636F1383EF238363239383EF2393231383376F138303),
    .INIT_08(256'h2323136713671367136713671367138303833313EF1393133393B393EF139333),
    .INIT_09(256'hE71383671383038363931323B7372323136FE71383671383038363931323B737),
    .INIT_0A(256'hEFEFEF23136F13830313EF239313931393139313B7373723136F1383EF23136F),
    .INIT_0B(256'h83038363839393232323232323231367131383EF231367131383EFEFEFEFEFEF),
    .INIT_0C(256'h830313EFEF1363EF13E7136383EF2323232313038303631383EF671383038303),
    .INIT_0D(256'hEF239313931393139313B73713132337136FEF23136FEF13EF6F138303830383),
    .INIT_0E(256'hEF13EF13230313EF671313038303836383931323232323136713376F13830313),
    .INIT_0F(256'h8363038363836F23232323930367131303836393638303EF232323131323136F),
    .INIT_10(256'h2313671313830383A32323239383EF2313232393139323136F836F2323232313),
    .INIT_11(256'h8367130383038313EF23936383EF232323932323136713130383EF13EF231313),
    .INIT_12(256'h132323136F936F03EFEF13EF13EF139313936383EF1313930323EF136F13EF63),
    .INIT_13(256'h93232323231363936F13239383671313830383EF63EF1313EF1363930393EF23),
    .INIT_14(256'h938303EF23231323239313932313671367131303830383EFEF2313EF1313EF13),
    .INIT_15(256'h136713130383EF13EF13EF23131323136713138303832323232323A323932323),
    .INIT_16(256'h038303830383038313EF63836313938303EF93EF232323132323232313232323),
    .INIT_17(256'h63939383EFE303EFEF13EF13EF13931313EF6383EF1393036F13632383671383),
    .INIT_18(256'h13EFEF13EF1363132313032363932393B393938383E3030313236333B3B383EF),
    .INIT_19(256'h639383EF93EF232323232313132323232323136F136FEF136F236F93136F236F),
    .INIT_1A(256'h13EF6383EF1393036F2393EF13632383671383038303830383038313EF631383),
    .INIT_1B(256'h9383B3138383E30313236333B3B383EF63939383EFE303EFEF13EF13EF139313),
    .INIT_1C(256'h231363936FEF136F9313136F236F13EFEF13EF13631323130323632393832393),
    .INIT_1D(256'h6F132393938383EF23136713671313830383EFEF232313EF13EF1393EF132323),
    .INIT_1E(256'h1393639313932323232323232323B7132323231367036F132393938383EF2313),
    .INIT_1F(256'h830383EF13931303EF23232323231393639393939333636393E313936F131363),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_008,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  // address_offset=2048;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00005328A08A513C48157E3DFE52E87FEC030710F31A5F3FFFE10018403959E3),
    .INITP_01(256'hEA20280181000000143467402050C2401000100460050C09800C6003000000E0),
    .INITP_02(256'h08944CA00068400000A0000000100092809004020A40080B00B40008000004EA),
    .INITP_03(256'h0802820100020264990011480D14812BF29108944C94000C900016A5204FE491),
    .INIT_00(256'h03F808C2636B12460882F8C3AB130802A2C2BAEBEA8E03F88EC3AB130882C6EB),
    .INIT_01(256'hCECDAB2B0B038B83EB81EB4C034303F84E4DAA8A10421208028243F8F8428B42),
    .INIT_02(256'hF8C1C3EB130842F8420882E3EB13EA1308C2C2EA81C3EB821308C2C2038282B9),
    .INIT_03(256'hEBCDBA03EBF84E4D104202031208F8F882AA1208C2C3FBE3138B03F848034303),
    .INIT_04(256'hCEAB438B83EBEB1367EB13EA1308C2C2C385BBE381C3EB1208C283C2020239EB),
    .INIT_05(256'h4081B2BAA28BBA1340BAAAD213F8080242C2FBE381C3F8420882F8CECD7D03CD),
    .INIT_06(256'hD70BF08293928040D20B4040D30BD40B40D50BD60B40BAD2134081F3FBA3BA13),
    .INIT_07(256'h0A028A10829192930280A6108090089093CC90C3930897C39380930BF0809092),
    .INIT_08(256'h919280400240024002400240024080929290820A1082028AC2CBC38B10420202),
    .INIT_09(256'hC002134080929290364202932A2A919280F8C002134080929290364202932A2A),
    .INIT_0A(256'h08F0F0938008809092020893C2030383030404022A130B9280108090F89380F8),
    .INIT_0B(256'h929290CA130504929496979193958040800290F8938040800290080010F80810),
    .INIT_0C(256'h9092020808828E0882C082C313081011D09104131312C58513F0408095959494),
    .INIT_0D(256'h0893C2030383030404022A130282920B80F8F89380F8F00208F0809595949492),
    .INIT_0E(256'hF0820882971284F04080029492929008130282909391928040820A0880909202),
    .INIT_0F(256'hD378E3E3C413F8D511D690C3134080029290050300929308979293C2829680F8),
    .INIT_10(256'h92804080029292900215160F0393089382979602C3029580F8D3F8D5D1D650C3),
    .INIT_11(256'h9340809492929002F04FC3C36BF09394968297958040800292900802F8938282),
    .INIT_12(256'h82919280F802F81208F082084208420283022893F842828263940884F802F0CC),
    .INIT_13(256'h029091929380CF03F8020FC32B4080029292900802F04202088286031282F093),
    .INIT_14(256'h03939308929382979602C302958040024080029492929008F00F82F80284F082),
    .INIT_15(256'h8040800292900802F802F8938282928040800292929012131108080217031516),
    .INIT_16(256'h959595949492929002F0CE938804822B2BF08408979091C59392939482959697),
    .INIT_17(256'h28858293F08ED208F04208420842028384F82993F882C223F842CBD493408095),
    .INIT_18(256'h0208F0420882870208831209FBEB50CB43C3CA132B812B2BC493A4C2838593F8),
    .INIT_19(256'hCE822BF084089790919493C582929395969780F803F8F042F809F8C505F893F8),
    .INIT_1A(256'h84F82993F882C223F8D403F042CED493408095959595949492929002F0CC0493),
    .INIT_1B(256'hC35343CB132B872BC493A6C2838593F828858293F08BD208F042084208420283),
    .INIT_1C(256'h9380CF03F8F042F8C50504F893F80208F0420882860208831209F209EB2B10CB),
    .INIT_1D(256'hF08001FBC39023F09380400240800292929008F0110842F802F80282F0829192),
    .INIT_1E(256'h3DC4CAC4823A95969790919295972CC4939496804022F08001FBC39023F09380),
    .INIT_1F(256'h939393080202859308939495969702024B050285060328C03AC4063A00063C84),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_017,inst_doa_i2_016,inst_doa_i2_015,inst_doa_i2_014,inst_doa_i2_013,inst_doa_i2_012,inst_doa_i2_011,inst_doa_i2_010,inst_doa_i2_009}));
  // address_offset=2048;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h10E33A60828A5089110800BF877A0381DB1A7898190F12C1C5A2CB085E2C3BFB),
    .INITP_01(256'h02000002310041500404CC80010822000002040B8C6110C30000C0002008060A),
    .INITP_02(256'h04A0080200C8500080A1000010050100068010401850480C00A4082040000180),
    .INITP_03(256'h10808142047CE4E9335020006C84910002200D0840304014840034110C080421),
    .INIT_00(256'h04670442BFE1200764322705E120C442952939D9E1390C77BDFDE120A43281E1),
    .INIT_01(256'hB9B1414141FD41FDD981E1B92039FCF7A9A94141B49520545301011707013D95),
    .INIT_02(256'h078139D9203492A7057432A5D920E120E42D95E18139D9722070292D399599B1),
    .INIT_03(256'hE181353CD95781815495004020B4476795D920144201059120BD0407B9283934),
    .INIT_04(256'hB541054105E1D920BDD920E120B4523D95010591A53DE1206029312D9995B9D9),
    .INIT_05(256'h00A93DF591050520000505912067C44201810591A539C7056432A78181B93CB9),
    .INIT_06(256'h2100D7010420C000710000002D002900002D0029000005912000BD29F9910520),
    .INIT_07(256'h0D2905D001242004A0C081404030F43DF1013DFD01143D0504C0710097403020),
    .INIT_08(256'h2420C0000000000000000000FC00401020302109E09DA009290D29057001A029),
    .INIT_09(256'h01110100401020302551410400002420C0770111010040102030254131040000),
    .INIT_0A(256'h50D3D704C0C4403020307404A11100010008503000000020C0644030C704C077),
    .INIT_0B(256'h506070CD50045050482004544C248000400030F704C000400030A4B05057E430),
    .INIT_0C(256'h706002347002D5B00201020171342121393DB10111504D015047008010203040),
    .INIT_0D(256'hD404C1B10001001C8001000001012000C0F74704C01737028467801020304050),
    .INIT_0E(256'hD70294B12501012700400000102030BD01FC0148042420C00001002440302001),
    .INIT_0F(256'h11B985D5210157213D393D51110080006070BD04812030A4042C3001012080F7),
    .INIT_10(256'h20C0008000506070353D3D255130803401042008010124804701973D39353951),
    .INIT_11(256'h3000804050607000533DFD8171832C4820010424800040002030D00157045101),
    .INIT_12(256'h012420C0070007C1706302F401F401003011BC30675101012581640167F8B301),
    .INIT_13(256'h0148242004C03D0427003D05710040001020302001230104F4B1BD5151019304),
    .INIT_14(256'h513020D03834010420140101248000FC00400000102030605325024751019301),
    .INIT_15(256'h000040002030900117A13704510120C0008000506070BDBD8181B53925A13D3D),
    .INIT_16(256'h8090A0B0C0D0E0F0F46381303D00018189C301F05CD8D40130D0CCC801A4A084),
    .INIT_17(256'hBC020130F381C2605301E402E40200300183BC3067020225F701018230000070),
    .INIT_18(256'h0000F301B4B1A151B90551BD314151412D05097191B18189022881293E493063),
    .INIT_19(256'h010189E301105CD8D4C8300101D0CCA4A084003700573301E7813712A1570087),
    .INIT_1A(256'h0183BC3067020225D7BEF883010182300000708090A0B0C0D0E0F0F893010030),
    .INIT_1B(256'h0501310971990189022881293E493063BC020130F381C2605301E402E4020030),
    .INIT_1C(256'h04C03D046723010712510037003700E0D30190B1A1A1B9FDA18135BD41813641),
    .INIT_1D(256'hD3403CFD0530102304C000FC004000102030100381810107A127510173012420),
    .INIT_1E(256'h425201E20102E4E0DC585450240400014C482080001033403CFDFD30108304C0),
    .INIT_1F(256'h605040F401280130643034383C4001285D280080B43001810A81C0064080FA02),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_026,inst_doa_i2_025,inst_doa_i2_024,inst_doa_i2_023,inst_doa_i2_022,inst_doa_i2_021,inst_doa_i2_020,inst_doa_i2_019,inst_doa_i2_018}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h04103345A00C6DB0420A8BE2B4588220A2C59988881408942148A10028800248),
    .INITP_01(256'hAA294579200085333108898EA002AC4601904AB52B4D5F5424BC929CB55469A7),
    .INITP_02(256'hF674406020800A20050011162BAB0412124463D4116400040000A511A40051B8),
    .INITP_03(256'h85503DB0893A7E4C5AF988A6AE23014902DA0604580CA9241296B1EFB7DD88E4),
    .INIT_00(256'h6F133313136363633313936393932393E393B3936393936FE3A3939383331303),
    .INIT_01(256'h13E3B31323636F93B313631313236363333313136313E3B31323636F13136F93),
    .INIT_02(256'h9323636F1323033313636F93339363639393E3331323636F33136F3333131363),
    .INIT_03(256'h136F03E3EF67138303B763EF231367133383038303830383038303831363E3B3),
    .INIT_04(256'h936393136F13E3EF671383133763EF23136F23E3EF6713038323B763EF132323),
    .INIT_05(256'h23932323236FB3931363B3133313B3939363339393B33313B313936763339363),
    .INIT_06(256'hB39313E33323032303230323139303676313936393B36393136FA3936F23136F),
    .INIT_07(256'h63B3636F2313B303B36F23133383336F93B313936F33B3B393136333931333B3),
    .INIT_08(256'h13E3B3138383B3B36F9363136F9367E323933383336F23333303336763939393),
    .INIT_09(256'h136FA36763933363A39393039393636733E36313631393631313839383131367),
    .INIT_0A(256'h63633383936F93136733636303836713E313639393B383B383B36F93631367E3),
    .INIT_0B(256'h6F1363333393EF131363EF932323232323131323136F9367336303936F936713),
    .INIT_0C(256'h9313B32323232323232323232323132313671303830383038313E3EF93139313),
    .INIT_0D(256'h8303830383038333236363E38313139313236363136F139313931337B7931363),
    .INIT_0E(256'h6393136F13636F13636F13636F13E393831313636F1393131367130383038303),
    .INIT_0F(256'h33E3939303E313936F9393631313938363939303E393831393331333936F1313),
    .INIT_10(256'h832393636393636393636393039363139303939363E393039313B393B3936F13),
    .INIT_11(256'h93E39363936363936F9313E39363936F136F93936F93138363936F13A3636313),
    .INIT_12(256'h636F939363136F93EF139333639303E313E39313E39393E3936F039393131363),
    .INIT_13(256'h23232313936313836F1323636F9363B3133313238363931333136393E3931323),
    .INIT_14(256'h336F9363B31333339363936393E313931323636F1393631393636303039383EF),
    .INIT_15(256'h2323239323136FA36F13136F936F936F93136F1323636F1323636F932383B363),
    .INIT_16(256'h372313676F6367671383EF232323232323231323136F931393671383EF232323),
    .INIT_17(256'h13133737EF1337EF2313133767130383EF13EF23232323232313939313232323),
    .INIT_18(256'h1363B3B767130333131363B393B7671303B3639313B7636F13133783EF931393),
    .INIT_19(256'h232323131323136713E39313673313638313931393676713033313671303B393),
    .INIT_1A(256'h6F13038303830323232323839303EFEF1313932393EF639383EF13EF13932323),
    .INIT_1B(256'h632323232323136713036713036F13032323232383930383EF13232323136F83),
    .INIT_1C(256'hB76F036713830383038313EF63EF139313136F13EF639303EF03EF2393631313),
    .INIT_1D(256'h23136F13132313830333139313EF2313036723239323232313E3932323139323),
    .INIT_1E(256'h136FEF6F13830313EF6393139323832363130383B3931393EF03631383B7EF23),
    .INIT_1F(256'h03EF132323136F1323B3038383232323238303B39313239393930383EF132323),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_008,inst_doa_i3_007,inst_doa_i3_006,inst_doa_i3_005,inst_doa_i3_004,inst_doa_i3_003,inst_doa_i3_002,inst_doa_i3_001,inst_doa_i3_000}));
  // address_offset=3072;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h1F590DF277FE9A7FFFADC3CD4802404840900005F30211359C28ACFE08A080E8),
    .INITP_01(256'h54188D78B6DB90000019121180000010122006EDF471FE89EFE2FFC0FC29D6E5),
    .INITP_02(256'hBB10A0000820048803F52239587704C1088D019412B00901561558A20B6229FE),
    .INITP_03(256'h4242B58870C81CAA2004107D400400840004308280232018007680465328F528),
    .INIT_00(256'h00040203832A4308833CC36A430280030D4E1E3ECC063A000847454222C58394),
    .INIT_01(256'h83248203003A00020302810283003A4583028303AA83248203003AF82B3DF806),
    .INIT_02(256'hC3C0FAF88280230383BD00028383CD42420364438280BAF80203F883028303AA),
    .INIT_03(256'h80F8928208408090D20B86F89380408082969695959595949492929003AA2403),
    .INIT_04(256'hBBBC8303F8828208408090820A86F89380F894810840809290D00B87F8829392),
    .INIT_05(256'hD7C3D2D1D0F8C37B7B338404C1C3833B3B7544038384B3CBB3CBFB40C9C383C5),
    .INIT_06(256'h838B2B754497D496D495D49483C3D440880383C0FBB3BD8303F8C7C3F81703F8),
    .INIT_07(256'hBBC3FDF84083C364C3F81083C414C4F803C483C3F803C2C38B2B6404030303C2),
    .INIT_08(256'hC2C7C38363E3C38300030B03F803400B80C383A3C3F88083C3A44340CAC30322),
    .INIT_09(256'h43F8C740CAC3C38FC703C3E3C2830040C2CCCA433244C33243C4E3C2A3820340),
    .INIT_0A(256'hB342C3E383F8C28240C2C3C2E3A340C24C83CBEBCB43E3C3E38300030B03404B),
    .INIT_0B(256'h00026B020582F8028480F8C49294959793C2829680F8C340C28BE383F8C34082),
    .INIT_0C(256'h4286859495909192939596979697C494804080959494929290028FF84202C283),
    .INIT_0D(256'h9595949492929002003A83CF2382430202003AC3030005C40505022D8405A4FB),
    .INIT_0E(256'h7103C3F834CBF834CBF834CBF834CB02234334C8000203030440809696969595),
    .INIT_0F(256'h03AEC202D3CA030300040372C24303630F0303633843638342838BC38B000303),
    .INIT_10(256'h6300033B070370060372000363420EBB03620203EA788322C303C3CB43CBF834),
    .INIT_11(256'h030E03070375070300033408030003F802F80302F8C243D3CD03F80200BAC002),
    .INIT_12(256'h3A0003830E3CF842F802C23BCA3AD38D0387C603090304060300D303C603348B),
    .INIT_13(256'h91929342064AC6D6F88280BAF8C2238303030200D33BC383C303228324C30200),
    .INIT_14(256'h03F8826283038302036A43E30363838302003A0003830A3CC3EA2B93948393F8),
    .INIT_15(256'h959497839380F8C7F82B0BF803F842F80334F802003AF88280BAF8C300E2423C),
    .INIT_16(256'h0A968040E08240408090F893979695949397839280F802C303408090F8939796),
    .INIT_17(256'h83822A2BF8822AF89382802A40809290E002F893979695949702028383939291),
    .INIT_18(256'hAAC7BB834082A243BBAAC7BBC383408262438543BB2B80F880822A90F8020303),
    .INIT_19(256'h949597C2829680400289438340C28ACC5203030303404082A242AA4082E243BB),
    .INIT_1A(256'hE880959494929214911391900393E8F802030202F4004F83920084F805C49293),
    .INIT_1B(256'h8597909192938040BAA240AA82E880921314905190031313E88282939280F852),
    .INIT_1C(256'h0BF8944080949492929002008AF802C203820002008C8294F892009384B30203),
    .INIT_1D(256'h9280E0808213839092828A0382F89380124015D10314130203CDC3D0D1C303C9),
    .INIT_1E(256'h80F8E0E880909202E8CFC282FB02231381C312D2C34B0383F812CB82CB0BE893),
    .INIT_1F(256'h13E082939280E08014F392131315D1169090D3C3038B05F3FB032323E8829392),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_017,inst_doa_i3_016,inst_doa_i3_015,inst_doa_i3_014,inst_doa_i3_013,inst_doa_i3_012,inst_doa_i3_011,inst_doa_i3_010,inst_doa_i3_009}));
  // address_offset=3072;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hB000000017F0006C800080200B12D040D8950FF21000E1244228221009008040),
    .INITP_01(256'h0698CD00B24A0020001013060000803800400C080400800160D2402840090405),
    .INITP_02(256'h0464002020A00A2007974200400600000088001C0281DA80FB8A000203938680),
    .INITP_03(256'h06000880F00A4328421D00470004482402840004000206000240000100800948),
    .INIT_00(256'h90803901FD3803823546013D0104B4C08117642201AC12B081AE060502520170),
    .INIT_01(256'h01AC3105614930C035010205FD6549033131FD000101AC31054149E7113DE700),
    .INIT_02(256'h052D4937053101258049B08039010135FDFCB129052D49573901173131FD0001),
    .INIT_03(256'hC0A7C181000040308100016704C0008039D0E0F000102030405060700001B43D),
    .INIT_04(256'h0D31010CA7C181300040308100019704C097A1810000402030A1000177010420),
    .INIT_05(256'hB9413939398735310DC6300C35013D3DC1C13E3C01313D413D21FD0031310101),
    .INIT_06(256'h351111413EC1F1C1E1C1D1C141410100B10001010D2D31013CD7AD0527B911D7),
    .INIT_07(256'h353129374105390139E74611390239B73C310101373535350909C1390C003535),
    .INIT_08(256'h010135050101393980003900D70000BD35053D013D87413931013D003DFD00FD),
    .INIT_09(256'h01C7810031053101B9FD05FD050101003901398141FD814101FDFD05FD056400),
    .INIT_0A(256'h2D01290101870505003939010101000101050161613D01390139B00039000001),
    .INIT_0B(256'h700049262901B7010101F701504824044C01012080B705002901010197050001),
    .INIT_0C(256'h0101496864D8D4D0CCA4A084605C01C8000080203040506070010107FD010202),
    .INIT_0D(256'h90A0B0C0D0E0F061015D020101010501053D5DB9949082FE80AC030000FCFD2A),
    .INIT_0E(256'hB92441270629578235872259B742B905050112D540C08CB40000004050607080),
    .INIT_0F(256'h388111090135FCA81024002941052405B5FCB801BD4101410535053909702400),
    .INIT_10(256'h013D945DBD94B135603135A40105B5EDA001010001B64101410529053D09B742),
    .INIT_11(256'hFCB5C035BCB1B5CC50280AB590B58C37000700010711090135A8C7093D5D0105),
    .INIT_12(256'h5D408001824287035301024D010A0131A03111B04540E0B5D4F0014011200635),
    .INIT_13(256'h40383C03020311019705315DE701342980390535015D1105390438FDBCFD0535),
    .INIT_14(256'h3D3703BD2980393D000101B500BDFD0105315D508001824201293C2010013047),
    .INIT_15(256'hBCB804B0B400F782E741418720F7FDC740024705315D2705315DF7052D013F5D),
    .INIT_16(256'h002000003701000000702730C4C0BCB8B404A0B00057FC0101000070C734C4C0),
    .INIT_17(256'h6191000027D1005704A1C00000006070F7E12734C4C0BCB804E1FC9001B4B0AC),
    .INIT_18(256'h41013D3F0025A139FD21013D01000005A13901E1FD00015740110030A70C040C),
    .INIT_19(256'h482404010120800000B14105002911290110000000000065A129610045A13DFD),
    .INIT_1A(256'hD3802030405060253E393D70311293130120024D02503D1212F001770101504C),
    .INIT_1B(256'h814CC8A4A0844000FD21007D21A340203D3D3539303141313301010420C08701),
    .INIT_1C(256'h00C70200C0708090A0B001B08103010220D28000402611114730002C012D0030),
    .INIT_1D(256'h20C057402138B130013D0D20FD7704C040003C3D500000381CB9213D3D012081),
    .INIT_1E(256'hC0A777034030200173012171FD341038B9B13001390D20FD2740010191009304),
    .INIT_1F(256'h61C7010420C037403C3520E1403D353935301139200DBD05C151D5D173010420),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_026,inst_doa_i3_025,inst_doa_i3_024,inst_doa_i3_023,inst_doa_i3_022,inst_doa_i3_021,inst_doa_i3_020,inst_doa_i3_019,inst_doa_i3_018}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hD05CB00A04C90918AAA52B0700601D600C0114118248555502D2487CAB28D7C2),
    .INITP_01(256'h740B0A814016808832B12601A0150DE10D3205311656150605D13832B180AC29),
    .INITP_02(256'hB0C4014D072395D5412A81A0301AF279AABB051801325AA2A1D40B44C18014CC),
    .INITP_03(256'hB5A97A3766B2B25C1456A1027CACC8B321AC8C7035458DCFA798C05466640200),
    .INIT_00(256'h136F132393838337EF23136F13830323B39383836303B3931383232323239383),
    .INIT_01(256'h93EF23230323136703B76713836F13836F13836383EF2363239393938337EF23),
    .INIT_02(256'h1383036F232393232313836F13838303EF13EF1363836393EF13EF132393EF13),
    .INIT_03(256'h232313838303EF232323231323232393139323136F1383EF2323231323232313),
    .INIT_04(256'h9323232323232323A3132323378303EF9333B79303830383EF93131323232323),
    .INIT_05(256'h1363836393EF132393EF13EF639313832323136703671313830383EF13139393),
    .INIT_06(256'h93032323630303631303931383EF23136FEF23239323231383EF6713130383EF),
    .INIT_07(256'h93139383EF1323232313639313836FEF1367131383EFEF232323230333231313),
    .INIT_08(256'h13EF13931393EF131303EF2323232323136713671313830383EF13EF13EF2393),
    .INIT_09(256'hEF1323232313639313836F1383EF23136F6713130383038323639303EFEF13EF),
    .INIT_0A(256'hEF23A3132333138323136713671313830383EF13EF13EF132323232393930383),
    .INIT_0B(256'hEF23A3B31383EF136393939383EF132323232313231363936367131383EF6383),
    .INIT_0C(256'h83EF13EF6313232323232383231367136F6F23A3B3036713138303830383EF13),
    .INIT_0D(256'h23239303836F83671303830383038313EF638363EF139313136F13EF63036313),
    .INIT_0E(256'h671383038323232323232393A393038383EF2323231323239313932313672323),
    .INIT_0F(256'hA3931383EF1393EF1323232313671313830383EF13EF13EF1393EF1323232313),
    .INIT_10(256'h1313830383EFA3938323232323932393833763031393370313B7EF233383EFEF),
    .INIT_11(256'h136713830383A3931383EF13EF1393EF13232323136393836F93E3B363838367),
    .INIT_12(256'h23232323232323136FA393836F23836F23836F9383E393639367136363639367),
    .INIT_13(256'h83EF13E33313036F1383138303038303838303630393931393B7EF3793EF2323),
    .INIT_14(256'h93631393136363676723239337670363139303B76FEF13E3A393139383EFE703),
    .INIT_15(256'h6713EF6363936733EF93B36FB363336713EF9367E3139333B36313E393136363),
    .INIT_16(256'h6313936F93A393938363939367E3A393938363936393633393B36733EF33E3B3),
    .INIT_17(256'h9363131367E3E3239393036F2393232323232323230323938303038303838383),
    .INIT_18(256'hA323A323A323A323A323A323A32367B39793B36763E31323232323B313936363),
    .INIT_19(256'h936F9367E3A3930393639303936FE333339393E793B397936FB393B393936723),
    .INIT_1A(256'h2323131367136733E31363638383B3B3131363671333E303939367E3A3939303),
    .INIT_1B(256'h1393B73793EFEF1337EF13EF13931393B7B7EF2313931393231393B72313EF23),
    .INIT_1C(256'h6176726D76726FEF13EF13EF1393139313931393B73793EF13EF139313931393),
    .INIT_1D(256'h6155327431740D6F33636F68005F75006C7320752E6920610D0D742E6920610D),
    .INIT_1E(256'h73645F006C5F6C6F6173645F655F6C006973645F002E64730021726F20726E65),
    .INIT_1F(256'h6D2D255F0A696F6E2D2F250A652D6F486E72645F655F6C646873645F005F6C65),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i4_008,inst_doa_i4_007,inst_doa_i4_006,inst_doa_i4_005,inst_doa_i4_004,inst_doa_i4_003,inst_doa_i4_002,inst_doa_i4_001,inst_doa_i4_000}));
  // address_offset=4096;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h883387FDFFC4C441441C00080009F0B0020049281110A882408496FA5A90CF0C),
    .INITP_01(256'h4900152000044020C400CA105800C80282060006840028308324804C02200045),
    .INITP_02(256'hC75FFA00FD468AA8A2914E1D40736F666120002400AB9008012906FA052B9DAB),
    .INITP_03(256'h20823252AA5256101446A51A37520D4836D1F09201FC679A6E77F581FFFF6FFD),
    .INIT_00(256'h80E08089C390AB0BE09380E080909214FBE313138ED3C3CB0323161590510313),
    .INIT_01(256'h82E0919312928040EA0B408090E08090F88090C713E0892089EBCBC3AB0BE093),
    .INIT_02(256'h809393F816150351150313F880929092E042F802CA138C03F80200020503F802),
    .INIT_03(256'h161203939393F8959697938294929302C3029180F88090F89596508311949303),
    .INIT_04(256'h031514051410171605020517239494E0430323C312121313F80282C313111015),
    .INIT_05(256'h02C8138A03F80205030002F8C2FB82A393928040124080029292900003030302),
    .INIT_06(256'hC3E3901104D3D38FBBE3830313E09380F8E016150351150313E04080029290F8),
    .INIT_07(256'hFB028223E08291929380C8FB03A3F8E04240800290F8E0D591D6109383D6030B),
    .INIT_08(256'h420042028302F8028412E09394959697804002408002929290E0420002F805F3),
    .INIT_09(256'hE08291929380CBFB03A3F88090E89380F840800294929290148A0313F8E08200),
    .INIT_0A(256'hF8858503968B03A393804002408002929290F802E04200021516905182031313),
    .INIT_0B(256'hF816054A02A3F8024B7A840322E00497939495829680CF03C040800290F8C213),
    .INIT_0C(256'h94F802F8C28593949697921395804002F8F81605CBA34080029494929290E0C2),
    .INIT_0D(256'h9051839393F8D4408095949492929002F8C2138DF0020203C20002F80512CE84),
    .INIT_0E(256'h40809292901516111210170302FB939393F891929382979602C3029580409596),
    .INIT_0F(256'h02FB4223F80282E08291929380408002929290F802E042F80282E08291929380),
    .INIT_10(256'h8002929290E002F32316D01591031243130B0CD323C30394C30BE012C213E8E0),
    .INIT_11(256'h02408092929002FB0223E042F80282E08291929380C5FBA3F883394343129340),
    .INIT_12(256'h9394959790919380F882FBA3F89113F8109300F3A3CB03C4034002C5E4C40340),
    .INIT_13(256'h13F80271C20512E080954295959594949290920D920562858502E00C84E89692),
    .INIT_14(256'h03060282C3E3A0404093D1830B40928202C3D30BF8F8028B05FBFB8423E8C012),
    .INIT_15(256'h40C2F8A6E5414002F84102F802EC0240C2F841404B2B6BB2C2F302354B0B2C3D),
    .INIT_16(256'hFA43BBF8FBC7C2C3E34783BB40F4C7C2C3E3BE83F103CB83FBE34002F802AC02),
    .INIT_17(256'hBBBF830140F4F4D7C2C3D3F8D7C3D7D6D5D4D3D2D1D4D0C2D4D1D7D7D7D7D1D1),
    .INIT_18(256'h80808081818181828282828383834043014B83400AB38393929190433B3BC9C8),
    .INIT_19(256'h83F843408CC7C3E3C28FC3E383F8BC0383C34040414301CBF8F2CBF2CBFA4080),
    .INIT_1A(256'h92930280400240C2C98383CC63E3C3830303054082C28EE3C383408CC7C2C3E3),
    .INIT_1B(256'h04042A0B02E0F0822AD802E002C203430A2BE8CA02C20303D103032A1002E091),
    .INIT_1C(256'h36AFB4322FB4F8F802F842F842C20303030304042A0B02F842F842C203030303),
    .INIT_1D(256'h37A700B000B0053919371032003430002FB4063A17B7B9B905059097B7B9B905),
    .INIT_1E(256'hBA2FAF00B1B6B43C34BA2FAF39BAB400B6BA2FAF0017B7B40090B9B1123ABA32),
    .INIT_1F(256'hB000392F0039373116003900302A103200B92FAF303AB400B9BA2FAF00B9B436),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_004096_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i4_017,inst_doa_i4_016,inst_doa_i4_015,inst_doa_i4_014,inst_doa_i4_013,inst_doa_i4_012,inst_doa_i4_011,inst_doa_i4_010,inst_doa_i4_009}));
  // address_offset=4096;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h806304020905C0002420201864419080000019019000A4320284029892B04080),
    .INITP_01(256'h410811010004000800008890100440000084040480502300062100290620A00C),
    .INITP_02(256'h07080400F406000A200008102650E0CC55000B040129040081210C000402AC82),
    .INITP_03(256'h828372562256533481D24E9D039410104501202810804B184D02408400000404),
    .INIT_00(256'hC0E740BD053091003704C0874030203C35FD40E13D01390D20D53D3D35395151),
    .INIT_01(256'h01C724043020C0009100004030A74030F7403001302781BCBD4141FD91009704),
    .INIT_02(256'hC06151273D355039385150A740103020D701570181C1BD04C701B011BD109701),
    .INIT_03(256'h31B951705060073C3834440140A084040101A440374030773939315135B904F8),
    .INIT_04(256'h018181818145C581C111C12900304027913D00F18191A1B1538C0101BDB5A531),
    .INIT_05(256'h0181C1BD049701BD10A01167013D01D10420C0003000C00090A0B0F0D1000001),
    .INIT_06(256'h51D53139396151313DD10104308704C027E73D35503938515047004000203027),
    .INIT_07(256'hC10101D1F701242004C0B93D04D1A7C70100400030473739353135113135200D),
    .INIT_08(256'h013001003011970101305728482420048000FC0040001020306701401187BD09),
    .INIT_09(256'hB701242004C0B93D08D1A740303704C00700800040506070813DF8C1B7A70230),
    .INIT_0A(256'h77B9B508B93504D904C000FC00400010203027011701F0113D3D353901516151),
    .INIT_0B(256'h07A5BD3D010217013D3D0104D18701044C48240120803D088100400030C70130),
    .INIT_0C(256'h11D3049701014C4820045030248000007727BDB939020080003040506070B702),
    .INIT_0D(256'h353951615177020080203040506070010701308177010220D2A000B781304A11),
    .INIT_0E(256'h00805060703D3DB981B525513DF9203010B33C38340104202801012480003D3D),
    .INIT_0F(256'h3DF901250701012301242004C0004000102030630127013701015701242004C0),
    .INIT_10(256'h4000102030233D05253D35393551B505A1003E01F9B10011B10053A9299157C3),
    .INIT_11(256'hFC00401020303DF900257301870101A301242004C00105255701B52D2DA15100),
    .INIT_12(256'h5C58544CC8A48440E73DF52527BD01573D91900925BD0CBD080000812DBD0400),
    .INIT_13(256'h21D702292AB15143C05002304060708090B0A0D9B20CF9B201005300014750A0),
    .INIT_14(256'h0481FC010181810000BD3DB10000513DFCB1B1000797025DBDF90D01D5470131),
    .INIT_15(256'h0001E7010100002847002C772C01280001D7000081050535313100AD0505302D),
    .INIT_16(256'hB181F1A70DB505050101010D00B9B5050501B901B10C01310D29002C8728812C),
    .INIT_17(256'h3DB0013C0039B5B1111101B7C19145197175797D15F11D917161514131211101),
    .INIT_18(256'h2D2D2D2D2D2D2D2D2D2D2D2D2D2D31150009300001B5412D2D2D2D393DC10181),
    .INIT_19(256'h0167010081B905FD0501050101F7B03D3DC1008100150009B735413521FD002D),
    .INIT_1A(256'h200400C000000035810531350101393900FD8100FD2981FD05010081B9050501),
    .INIT_1B(256'h10900000C117474100E71003108100110000B73941E100000140000020803324),
    .INIT_1C(256'h1BD9DC1C5DDCE773D003018301C1F100A10010900000A1E3016301A16100C100),
    .INIT_1D(256'h190B00DC00DC001BC89C5C1B005C1C001C190288C8999D9A0800105B999D5A08),
    .INIT_1E(256'hD75B58001B581C009B575B58005A1C0099175B58008B9D1D00881958191C9948),
    .INIT_1F(256'h1A000200009D085D51000000599A141B00DA5D58199A1C0059175B5800591C00),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_004096_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i4_026,inst_doa_i4_025,inst_doa_i4_024,inst_doa_i4_023,inst_doa_i4_022,inst_doa_i4_021,inst_doa_i4_020,inst_doa_i4_019,inst_doa_i4_018}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h000000000039D4B145B57E41B777D0920132D37FF5678482BB1FFE14A597F573),
    .INITP_01(256'h00A595E7FA000A0036DB6DB6DB6DB6DB647B2443A5A57FD5561062F042000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h2572740A6420302A253A6420302A252D2D2D2D2D2D2000652070207374732562),
    .INIT_01(256'h6300747464647661202578782A252D2D2D2D2D2D2D2D200A6620746D20646573),
    .INIT_02(256'h2D202D2D2D2D20206F20696664202073612070207374697325617400303A7465),
    .INIT_03(256'h322038303020006E20007320007420007020006420332A25002D2D2D202D202D),
    .INIT_04(256'h5F00645F25302A2525302A25002D2D2D20200A72647320732565707333787820),
    .INIT_05(256'h006D00736C7464666E6163250A556E5773206D5425645F3A6163656468526C64),
    .INIT_06(256'h0203020402030200006338343000433834306574006D082008002525083E6866),
    .INIT_07(256'h0203020402030207020302040203020502030204020302060203020402030205),
    .INIT_08(256'h20202D007C0A4C28020302040203020502030204020302060203020402030205),
    .INIT_09(256'h0C30D0740A74652D796879203236200A64622E6420202030334A655369656468),
    .INIT_0A(256'h76006C002E552047147CB4702484B47CB4B05CA45C9090849074806480500C44),
    .INIT_0B(256'h040101C44A00017600696963672F2D692E2F2E000001FB0002655C6C646F6869),
    .INIT_0C(256'h0101040101040102040101040101040102040101040101040101040101040101),
    .INIT_0D(256'h0404010104010204010204010104010104010404010104010204010104010104),
    .INIT_0E(256'h2F626376722F2E2E0000B4640002021C00002503111100000000000001570001),
    .INIT_0F(256'h0031205563696C776E336965736C2D2D756C2F76696C2D2D696E652F76767266),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i5_008,inst_doa_i5_007,inst_doa_i5_006,inst_doa_i5_005,inst_doa_i5_004,inst_doa_i5_003,inst_doa_i5_002,inst_doa_i5_001,inst_doa_i5_000}));
  // address_offset=5120;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h000000000018C08112107210999003A80102810000E5C0A29006001480830052),
    .INITP_01(256'h2EB553FBDF1039F00002002000082080057BE0B9ABFFFFFFF090003A28000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h1600B40090121A39160090121A39161696969696109600303A32B934B9901637),
    .INIT_01(256'h3A003234B205303100181012391616969616969696969600B61010B210B4B910),
    .INIT_02(256'h96969696909690963932B13A10BAB634B190101010301010163234001C18B437),
    .INIT_03(256'hB2903CBC1C180034B90032310010340032B9003CB93239160096969696969696),
    .INIT_04(256'hAF002FAF321939163219391600969696969600B210B890101600B4B232901210),
    .INIT_05(256'h00390034363917B73737B73900B9B632903030B7392FAF0537B73690B9AA382F),
    .INIT_06(256'h808080808080808000B29C1A1800A29C1A18003400B010049200B93100001034),
    .INIT_07(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_08(256'h10161000901014A7808080808080808080808080808080808080808080808080),
    .INIT_09(256'h0A27082A00B2303A103AB9A19890190090BA1297102E1719183A36BCB7B990B9),
    .INIT_0A(256'h3200B400191494A10C290C29082A082A08270A270A270B270B27092709270A27),
    .INIT_0B(256'h800104800102009700B9B337B1B6B3B997171780008087800000121212003237),
    .INIT_0C(256'h8104808104808104808104800104808104800104808104800104808104808104),
    .INIT_0D(256'h0080810480810480810480810480010480810480810480810480010480810480),
    .INIT_0E(256'hB1B31796B4171797000000250000800000008787000000F7C8B08C32CC010111),
    .INIT_0F(256'h0097199080B1B3B73599B999BA34B7B334B2B119B731BA33B9B317B49717B4B4),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_005120_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i5_017,inst_doa_i5_016,inst_doa_i5_015,inst_doa_i5_014,inst_doa_i5_013,inst_doa_i5_012,inst_doa_i5_011,inst_doa_i5_010,inst_doa_i5_009}));
  // address_offset=5120;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000529400052142459333D6808590831AFF1D44A40205F692ADB6EC56),
    .INITP_01(256'h0BEE83B1870234060000000000000000045970022200000004A05A14A1000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h8A005B00090C19488A00090C19488A024B4B4B0B484B00999A1BDD5E1E998A1E),
    .INIT_01(256'h9C00995DD8005D5D000E0C0C088A024B4B484B4B0B4B4B00D808085B5D18DA08),
    .INIT_02(256'h4B4B4B4B4B4B4B4B029C1A085B5C185E1A1C08C8085DC89C8A005C009E5ED81D),
    .INIT_03(256'h490908091E5E00DB9D0008DB00085B001BDD00085908488A008B0B4B4B0B4B0B),
    .INIT_04(256'h5800DC580219488A0E19488A008B4B4B4B4B00181D995C1D8A009B5B02090C08),
    .INIT_05(256'h001A001C005A029D1D195B0E00991EC808DC5B1B08005800D95B1B1C590B005A),
    .INIT_06(256'h0000000000000000009998CDCC009190CDCC0019009A02001C00C900000000DB),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h080814008B170015000000000000000000000000000000000000000000000000),
    .INIT_09(256'h000000000058199A1C88DA1B4C0B0C00C91A19094808080C881B021C19181359),
    .INIT_0A(256'hDC001C000B089190000000000000000000000000000000000000000000000000),
    .INIT_0B(256'hC04101C0C000001459988B9BD89AD8988BCB8B80404003401100000000001B1B),
    .INIT_0C(256'h4101C04001C04101C04001C04001C04001C04001C04001C04001C04001C04001),
    .INIT_0D(256'h40404001C04001C04001C04001C04001C04001C04001C04001C04001C04001C0),
    .INIT_0E(256'h9BD85BD9DCCB8B8B000000000001C0000000448644846095959592929500C000),
    .INIT_0F(256'h000CCBD091D90B4BDB4B988BD858D9D81B8B5D4C8B5ADB5B988BDC5B1459DCD9),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_005120_018 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i5_026,inst_doa_i5_025,inst_doa_i5_024,inst_doa_i5_023,inst_doa_i5_022,inst_doa_i5_021,inst_doa_i5_020,inst_doa_i5_019,inst_doa_i5_018}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i6_008,inst_doa_i6_007,inst_doa_i6_006,inst_doa_i6_005,inst_doa_i6_004,inst_doa_i6_003,inst_doa_i6_002,inst_doa_i6_001,inst_doa_i6_000}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i7_008,inst_doa_i7_007,inst_doa_i7_006,inst_doa_i7_005,inst_doa_i7_004,inst_doa_i7_003,inst_doa_i7_002,inst_doa_i7_001,inst_doa_i7_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b0/B0_2 ),
    .i1(\inst_doa_mux_b0/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b1/B0_2 ),
    .i1(\inst_doa_mux_b1/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i1_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_1  (
    .i0(inst_doa_i2_010),
    .i1(inst_doa_i3_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_2  (
    .i0(inst_doa_i4_010),
    .i1(inst_doa_i5_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_2 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_3 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b10/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b10/B0_2 ),
    .i1(\inst_doa_mux_b10/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b10/B1_0 ),
    .i1(\inst_doa_mux_b10/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i1_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_1  (
    .i0(inst_doa_i2_011),
    .i1(inst_doa_i3_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_2  (
    .i0(inst_doa_i4_011),
    .i1(inst_doa_i5_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_2 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_3 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b11/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b11/B0_2 ),
    .i1(\inst_doa_mux_b11/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b11/B1_0 ),
    .i1(\inst_doa_mux_b11/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_0  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i1_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_1  (
    .i0(inst_doa_i2_012),
    .i1(inst_doa_i3_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_2  (
    .i0(inst_doa_i4_012),
    .i1(inst_doa_i5_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_2 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_3 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b12/B0_0 ),
    .i1(\inst_doa_mux_b12/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b12/B0_2 ),
    .i1(\inst_doa_mux_b12/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b12/B1_0 ),
    .i1(\inst_doa_mux_b12/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[12]));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_0  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i1_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_1  (
    .i0(inst_doa_i2_013),
    .i1(inst_doa_i3_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_2  (
    .i0(inst_doa_i4_013),
    .i1(inst_doa_i5_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_2 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_3 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b13/B0_0 ),
    .i1(\inst_doa_mux_b13/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b13/B0_2 ),
    .i1(\inst_doa_mux_b13/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b13/B1_0 ),
    .i1(\inst_doa_mux_b13/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[13]));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_0  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i1_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_1  (
    .i0(inst_doa_i2_014),
    .i1(inst_doa_i3_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_2  (
    .i0(inst_doa_i4_014),
    .i1(inst_doa_i5_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_2 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_3 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b14/B0_0 ),
    .i1(\inst_doa_mux_b14/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b14/B0_2 ),
    .i1(\inst_doa_mux_b14/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b14/B1_0 ),
    .i1(\inst_doa_mux_b14/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[14]));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_0  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i1_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_1  (
    .i0(inst_doa_i2_015),
    .i1(inst_doa_i3_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_2  (
    .i0(inst_doa_i4_015),
    .i1(inst_doa_i5_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_2 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_3 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b15/B0_0 ),
    .i1(\inst_doa_mux_b15/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b15/B0_2 ),
    .i1(\inst_doa_mux_b15/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b15/B1_0 ),
    .i1(\inst_doa_mux_b15/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[15]));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_0  (
    .i0(inst_doa_i0_016),
    .i1(inst_doa_i1_016),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_0 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_1  (
    .i0(inst_doa_i2_016),
    .i1(inst_doa_i3_016),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_1 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_2  (
    .i0(inst_doa_i4_016),
    .i1(inst_doa_i5_016),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_2 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_3 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b16/B0_0 ),
    .i1(\inst_doa_mux_b16/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b16/B1_0 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b16/B0_2 ),
    .i1(\inst_doa_mux_b16/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b16/B1_1 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b16/B1_0 ),
    .i1(\inst_doa_mux_b16/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[16]));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_0  (
    .i0(inst_doa_i0_017),
    .i1(inst_doa_i1_017),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_0 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_1  (
    .i0(inst_doa_i2_017),
    .i1(inst_doa_i3_017),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_1 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_2  (
    .i0(inst_doa_i4_017),
    .i1(inst_doa_i5_017),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_2 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_3 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b17/B0_0 ),
    .i1(\inst_doa_mux_b17/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b17/B1_0 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b17/B0_2 ),
    .i1(\inst_doa_mux_b17/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b17/B1_1 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b17/B1_0 ),
    .i1(\inst_doa_mux_b17/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[17]));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_0  (
    .i0(inst_doa_i0_018),
    .i1(inst_doa_i1_018),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_0 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_1  (
    .i0(inst_doa_i2_018),
    .i1(inst_doa_i3_018),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_1 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_2  (
    .i0(inst_doa_i4_018),
    .i1(inst_doa_i5_018),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_2 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_3 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b18/B0_0 ),
    .i1(\inst_doa_mux_b18/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b18/B1_0 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b18/B0_2 ),
    .i1(\inst_doa_mux_b18/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b18/B1_1 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b18/B1_0 ),
    .i1(\inst_doa_mux_b18/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[18]));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_0  (
    .i0(inst_doa_i0_019),
    .i1(inst_doa_i1_019),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_0 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_1  (
    .i0(inst_doa_i2_019),
    .i1(inst_doa_i3_019),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_1 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_2  (
    .i0(inst_doa_i4_019),
    .i1(inst_doa_i5_019),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_2 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_3 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b19/B0_0 ),
    .i1(\inst_doa_mux_b19/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b19/B1_0 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b19/B0_2 ),
    .i1(\inst_doa_mux_b19/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b19/B1_1 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b19/B1_0 ),
    .i1(\inst_doa_mux_b19/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[19]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b2/B0_2 ),
    .i1(\inst_doa_mux_b2/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(\inst_doa_mux_b2/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_0  (
    .i0(inst_doa_i0_020),
    .i1(inst_doa_i1_020),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_0 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_1  (
    .i0(inst_doa_i2_020),
    .i1(inst_doa_i3_020),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_1 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_2  (
    .i0(inst_doa_i4_020),
    .i1(inst_doa_i5_020),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_2 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_3 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b20/B0_0 ),
    .i1(\inst_doa_mux_b20/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b20/B1_0 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b20/B0_2 ),
    .i1(\inst_doa_mux_b20/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b20/B1_1 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b20/B1_0 ),
    .i1(\inst_doa_mux_b20/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[20]));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_0  (
    .i0(inst_doa_i0_021),
    .i1(inst_doa_i1_021),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_0 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_1  (
    .i0(inst_doa_i2_021),
    .i1(inst_doa_i3_021),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_1 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_2  (
    .i0(inst_doa_i4_021),
    .i1(inst_doa_i5_021),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_2 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_3 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b21/B0_0 ),
    .i1(\inst_doa_mux_b21/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b21/B1_0 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b21/B0_2 ),
    .i1(\inst_doa_mux_b21/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b21/B1_1 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b21/B1_0 ),
    .i1(\inst_doa_mux_b21/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[21]));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_0  (
    .i0(inst_doa_i0_022),
    .i1(inst_doa_i1_022),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_0 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_1  (
    .i0(inst_doa_i2_022),
    .i1(inst_doa_i3_022),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_1 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_2  (
    .i0(inst_doa_i4_022),
    .i1(inst_doa_i5_022),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_2 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_3 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b22/B0_0 ),
    .i1(\inst_doa_mux_b22/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b22/B1_0 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b22/B0_2 ),
    .i1(\inst_doa_mux_b22/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b22/B1_1 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b22/B1_0 ),
    .i1(\inst_doa_mux_b22/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[22]));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_0  (
    .i0(inst_doa_i0_023),
    .i1(inst_doa_i1_023),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_0 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_1  (
    .i0(inst_doa_i2_023),
    .i1(inst_doa_i3_023),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_1 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_2  (
    .i0(inst_doa_i4_023),
    .i1(inst_doa_i5_023),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_2 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_3 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b23/B0_0 ),
    .i1(\inst_doa_mux_b23/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b23/B1_0 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b23/B0_2 ),
    .i1(\inst_doa_mux_b23/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b23/B1_1 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b23/B1_0 ),
    .i1(\inst_doa_mux_b23/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[23]));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_0  (
    .i0(inst_doa_i0_024),
    .i1(inst_doa_i1_024),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_0 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_1  (
    .i0(inst_doa_i2_024),
    .i1(inst_doa_i3_024),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_1 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_2  (
    .i0(inst_doa_i4_024),
    .i1(inst_doa_i5_024),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_2 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b24/B0_3 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b24/B0_0 ),
    .i1(\inst_doa_mux_b24/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b24/B1_0 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b24/B0_2 ),
    .i1(\inst_doa_mux_b24/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b24/B1_1 ));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b24/B1_0 ),
    .i1(\inst_doa_mux_b24/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[24]));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_0  (
    .i0(inst_doa_i0_025),
    .i1(inst_doa_i1_025),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_0 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_1  (
    .i0(inst_doa_i2_025),
    .i1(inst_doa_i3_025),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_1 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_2  (
    .i0(inst_doa_i4_025),
    .i1(inst_doa_i5_025),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_2 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b25/B0_3 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b25/B0_0 ),
    .i1(\inst_doa_mux_b25/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b25/B1_0 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b25/B0_2 ),
    .i1(\inst_doa_mux_b25/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b25/B1_1 ));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b25/B1_0 ),
    .i1(\inst_doa_mux_b25/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[25]));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_0  (
    .i0(inst_doa_i0_026),
    .i1(inst_doa_i1_026),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_0 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_1  (
    .i0(inst_doa_i2_026),
    .i1(inst_doa_i3_026),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_1 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_2  (
    .i0(inst_doa_i4_026),
    .i1(inst_doa_i5_026),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_2 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b26/B0_3 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b26/B0_0 ),
    .i1(\inst_doa_mux_b26/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b26/B1_0 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b26/B0_2 ),
    .i1(\inst_doa_mux_b26/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b26/B1_1 ));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b26/B1_0 ),
    .i1(\inst_doa_mux_b26/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[26]));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_0  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_0 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_1  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_1 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_2  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_2 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_3  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i0_027),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b27/B0_3 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b27/B0_0 ),
    .i1(\inst_doa_mux_b27/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b27/B1_0 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b27/B0_2 ),
    .i1(\inst_doa_mux_b27/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b27/B1_1 ));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b27/B1_0 ),
    .i1(\inst_doa_mux_b27/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[27]));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_0  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_0 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_1  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_1 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_2  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_2 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_3  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i0_028),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b28/B0_3 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b28/B0_0 ),
    .i1(\inst_doa_mux_b28/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b28/B1_0 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b28/B0_2 ),
    .i1(\inst_doa_mux_b28/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b28/B1_1 ));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b28/B1_0 ),
    .i1(\inst_doa_mux_b28/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[28]));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_0  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_0 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_1  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_1 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_2  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_2 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_3  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i0_029),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b29/B0_3 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b29/B0_0 ),
    .i1(\inst_doa_mux_b29/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b29/B1_0 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b29/B0_2 ),
    .i1(\inst_doa_mux_b29/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b29/B1_1 ));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b29/B1_0 ),
    .i1(\inst_doa_mux_b29/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[29]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i5_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b3/B0_2 ),
    .i1(\inst_doa_mux_b3/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b3/B1_0 ),
    .i1(\inst_doa_mux_b3/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_0  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_0 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_1  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_1 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_2  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_2 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_3  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i0_030),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b30/B0_3 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b30/B0_0 ),
    .i1(\inst_doa_mux_b30/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b30/B1_0 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b30/B0_2 ),
    .i1(\inst_doa_mux_b30/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b30/B1_1 ));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b30/B1_0 ),
    .i1(\inst_doa_mux_b30/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[30]));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_0  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_0 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_1  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_1 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_2  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_2 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_3  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i0_031),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b31/B0_3 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b31/B0_0 ),
    .i1(\inst_doa_mux_b31/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b31/B1_0 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b31/B0_2 ),
    .i1(\inst_doa_mux_b31/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b31/B1_1 ));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b31/B1_0 ),
    .i1(\inst_doa_mux_b31/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[31]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i5_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b4/B0_2 ),
    .i1(\inst_doa_mux_b4/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b4/B1_0 ),
    .i1(\inst_doa_mux_b4/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i5_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b5/B0_2 ),
    .i1(\inst_doa_mux_b5/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b5/B1_0 ),
    .i1(\inst_doa_mux_b5/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i5_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b6/B0_2 ),
    .i1(\inst_doa_mux_b6/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b6/B1_0 ),
    .i1(\inst_doa_mux_b6/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i5_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b7/B0_2 ),
    .i1(\inst_doa_mux_b7/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b7/B1_0 ),
    .i1(\inst_doa_mux_b7/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i5_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b8/B0_2 ),
    .i1(\inst_doa_mux_b8/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b8/B1_0 ),
    .i1(\inst_doa_mux_b8/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i1_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_1  (
    .i0(inst_doa_i2_009),
    .i1(inst_doa_i3_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_2  (
    .i0(inst_doa_i4_009),
    .i1(inst_doa_i5_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_2 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_3 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b9/B0_0 ),
    .i1(\inst_doa_mux_b9/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b9/B0_2 ),
    .i1(\inst_doa_mux_b9/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b9/B1_0 ),
    .i1(\inst_doa_mux_b9/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[9]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

